VERSION 5.5 ;

NAMESCASESENSITIVE ON ;

DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

UNITS
    DATABASE MICRONS 100  ;
END UNITS

MANUFACTURINGGRID    0.010000 ;

MACRO XOR3SP8V1_0
    CLASS CORE ;
    FOREIGN XOR3SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.66 1.46 2.10 1.74 ;
        END
    END IN2
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 20.34  LAYER ME1  ;
        ANTENNADIFFAREA 9.57  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.84  LAYER ME1  ;
        ANTENNAMAXAREACAR 24.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.38 1.92 9.66 2.52 ;
        RECT  9.38 0.62 9.66 1.22 ;
        RECT  9.38 0.62 9.54 2.52 ;
        RECT  8.42 1.52 9.54 1.68 ;
        RECT  8.42 1.46 8.72 1.74 ;
        RECT  8.34 1.92 8.62 2.52 ;
        RECT  8.34 0.62 8.62 1.22 ;
        RECT  8.42 0.62 8.58 2.52 ;
        END
    END OUT
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.64 1.38 7.94 1.76 ;
        END
    END IN3
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.78 1.42 1.18 1.70 ;
        END
    END IN1
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 10.40 3.48 ;
        RECT  9.94 2.88 10.22 3.48 ;
        RECT  9.90 1.92 10.18 2.52 ;
        RECT  9.96 1.92 10.12 3.48 ;
        RECT  8.86 1.92 9.14 2.52 ;
        RECT  8.92 1.92 9.08 3.48 ;
        RECT  7.82 1.92 8.10 2.52 ;
        RECT  7.88 1.92 8.04 3.48 ;
        RECT  1.72 1.92 2.00 2.20 ;
        RECT  1.82 1.92 1.98 3.48 ;
        RECT  0.72 1.86 1.00 2.14 ;
        RECT  0.78 1.86 0.94 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 10.40 0.28 ;
        RECT  9.94 -0.28 10.22 0.32 ;
        RECT  9.90 0.62 10.18 1.22 ;
        RECT  9.96 -0.28 10.12 1.22 ;
        RECT  8.86 0.62 9.14 1.22 ;
        RECT  8.92 -0.28 9.08 1.22 ;
        RECT  7.82 0.62 8.10 1.22 ;
        RECT  7.88 -0.28 8.04 1.22 ;
        RECT  1.48 -0.28 1.76 0.58 ;
        RECT  0.72 0.78 1.00 1.06 ;
        RECT  0.78 -0.28 0.94 1.06 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.20 0.78 0.48 1.06 ;
        RECT  0.20 1.86 0.48 2.14 ;
        RECT  0.22 0.78 0.38 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  2.24 0.76 2.52 1.04 ;
        RECT  2.28 1.22 2.66 1.50 ;
        RECT  2.28 0.76 2.44 2.20 ;
        RECT  2.24 1.92 2.52 2.20 ;
        RECT  2.72 0.76 3.00 1.04 ;
        RECT  2.82 0.76 2.98 2.20 ;
        RECT  2.72 1.92 3.00 2.20 ;
        RECT  2.72 1.92 2.88 2.63 ;
        RECT  2.58 2.35 2.88 2.63 ;
        RECT  1.92 0.44 3.92 0.60 ;
        RECT  3.76 0.44 3.92 1.04 ;
        RECT  1.92 0.44 2.08 0.94 ;
        RECT  1.24 0.78 2.08 0.94 ;
        RECT  3.76 0.76 4.04 1.04 ;
        RECT  1.24 0.78 1.52 1.06 ;
        RECT  3.82 0.76 3.98 2.20 ;
        RECT  1.24 1.86 1.52 2.14 ;
        RECT  3.76 1.92 4.04 2.20 ;
        RECT  1.34 0.78 1.50 2.68 ;
        RECT  1.34 2.40 1.66 2.68 ;
        RECT  4.80 0.76 5.08 1.04 ;
        RECT  4.92 1.54 5.22 1.82 ;
        RECT  4.92 0.76 5.08 2.20 ;
        RECT  4.80 1.92 5.08 2.20 ;
        RECT  3.24 0.76 3.52 1.04 ;
        RECT  5.40 0.76 5.68 1.04 ;
        RECT  5.46 0.76 5.62 2.20 ;
        RECT  3.30 0.76 3.46 2.20 ;
        RECT  3.24 1.92 3.52 2.20 ;
        RECT  5.40 1.92 5.68 2.20 ;
        RECT  3.36 1.92 3.52 2.52 ;
        RECT  5.40 1.92 5.56 2.52 ;
        RECT  3.36 2.36 5.56 2.52 ;
        RECT  4.40 0.44 6.60 0.60 ;
        RECT  4.40 0.44 4.56 1.04 ;
        RECT  4.28 0.76 4.56 1.04 ;
        RECT  6.44 0.76 6.72 1.04 ;
        RECT  4.34 0.76 4.50 2.20 ;
        RECT  6.44 0.44 6.60 2.20 ;
        RECT  4.28 1.92 4.56 2.20 ;
        RECT  6.44 1.92 6.72 2.20 ;
        RECT  5.92 0.76 6.20 1.04 ;
        RECT  5.98 0.76 6.14 2.20 ;
        RECT  5.92 1.92 6.20 2.20 ;
        RECT  6.04 1.92 6.20 2.70 ;
        RECT  6.04 2.54 7.42 2.70 ;
        RECT  7.14 2.48 7.42 2.76 ;
        RECT  7.26 0.76 7.54 1.04 ;
        RECT  7.12 1.14 7.42 1.42 ;
        RECT  7.26 0.76 7.42 2.20 ;
        RECT  7.26 1.92 7.54 2.20 ;
    END
END XOR3SP8V1_0

MACRO XOR3SP4V1_0
    CLASS CORE ;
    FOREIGN XOR3SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.64 1.38 7.94 1.76 ;
        END
    END IN3
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 18.45  LAYER ME1  ;
        ANTENNADIFFAREA 7.88  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.56  LAYER ME1  ;
        ANTENNAMAXAREACAR 33.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.42 1.46 8.72 1.74 ;
        RECT  8.34 1.92 8.62 2.52 ;
        RECT  8.34 0.62 8.62 1.22 ;
        RECT  8.42 0.62 8.58 2.52 ;
        END
    END OUT
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.66 1.46 2.10 1.74 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.78 1.42 1.18 1.70 ;
        END
    END IN1
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 9.60 3.48 ;
        RECT  8.98 2.88 9.42 3.48 ;
        RECT  8.98 1.92 9.14 3.48 ;
        RECT  8.86 1.92 9.14 2.52 ;
        RECT  7.82 1.92 8.10 2.52 ;
        RECT  7.88 1.92 8.04 3.48 ;
        RECT  1.72 1.92 2.00 2.20 ;
        RECT  1.82 1.92 1.98 3.48 ;
        RECT  0.72 1.86 1.00 2.14 ;
        RECT  0.78 1.86 0.94 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 9.60 0.28 ;
        RECT  8.98 -0.28 9.42 0.32 ;
        RECT  8.86 0.62 9.14 1.22 ;
        RECT  8.98 -0.28 9.14 1.22 ;
        RECT  7.82 0.62 8.10 1.22 ;
        RECT  7.88 -0.28 8.04 1.22 ;
        RECT  1.48 -0.28 1.76 0.58 ;
        RECT  0.72 0.78 1.00 1.06 ;
        RECT  0.78 -0.28 0.94 1.06 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.20 0.78 0.48 1.06 ;
        RECT  0.20 1.86 0.48 2.14 ;
        RECT  0.22 0.78 0.38 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  2.24 0.76 2.52 1.04 ;
        RECT  2.28 1.22 2.66 1.50 ;
        RECT  2.28 0.76 2.44 2.20 ;
        RECT  2.24 1.92 2.52 2.20 ;
        RECT  2.72 0.76 3.00 1.04 ;
        RECT  2.82 0.76 2.98 2.20 ;
        RECT  2.72 1.92 3.00 2.20 ;
        RECT  2.72 1.92 2.88 2.63 ;
        RECT  2.58 2.35 2.88 2.63 ;
        RECT  1.92 0.44 3.92 0.60 ;
        RECT  3.76 0.44 3.92 1.04 ;
        RECT  1.92 0.44 2.08 0.94 ;
        RECT  1.24 0.78 2.08 0.94 ;
        RECT  3.76 0.76 4.04 1.04 ;
        RECT  1.24 0.78 1.52 1.06 ;
        RECT  3.82 0.76 3.98 2.20 ;
        RECT  1.24 1.86 1.52 2.14 ;
        RECT  3.76 1.92 4.04 2.20 ;
        RECT  1.34 0.78 1.50 2.68 ;
        RECT  1.34 2.40 1.66 2.68 ;
        RECT  4.80 0.76 5.08 1.04 ;
        RECT  4.92 1.54 5.22 1.82 ;
        RECT  4.92 0.76 5.08 2.20 ;
        RECT  4.80 1.92 5.08 2.20 ;
        RECT  3.24 0.76 3.52 1.04 ;
        RECT  5.40 0.76 5.68 1.04 ;
        RECT  5.46 0.76 5.62 2.20 ;
        RECT  3.30 0.76 3.46 2.20 ;
        RECT  3.24 1.92 3.52 2.20 ;
        RECT  5.40 1.92 5.68 2.20 ;
        RECT  3.36 1.92 3.52 2.52 ;
        RECT  5.40 1.92 5.56 2.52 ;
        RECT  3.36 2.36 5.56 2.52 ;
        RECT  4.40 0.44 6.60 0.60 ;
        RECT  4.40 0.44 4.56 1.04 ;
        RECT  4.28 0.76 4.56 1.04 ;
        RECT  6.44 0.76 6.72 1.04 ;
        RECT  4.34 0.76 4.50 2.20 ;
        RECT  6.44 0.44 6.60 2.20 ;
        RECT  4.28 1.92 4.56 2.20 ;
        RECT  6.44 1.92 6.72 2.20 ;
        RECT  5.92 0.76 6.20 1.04 ;
        RECT  5.98 0.76 6.14 2.20 ;
        RECT  5.92 1.92 6.20 2.20 ;
        RECT  6.04 1.92 6.20 2.70 ;
        RECT  6.04 2.54 7.42 2.70 ;
        RECT  7.14 2.48 7.42 2.76 ;
        RECT  7.26 0.76 7.54 1.04 ;
        RECT  7.12 1.14 7.42 1.42 ;
        RECT  7.26 0.76 7.42 2.20 ;
        RECT  7.26 1.92 7.54 2.20 ;
    END
END XOR3SP4V1_0

MACRO XOR3SP2V1_0
    CLASS CORE ;
    FOREIGN XOR3SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.66 1.46 2.10 1.74 ;
        END
    END IN2
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 17.10  LAYER ME1  ;
        ANTENNADIFFAREA 6.91  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.41  LAYER ME1  ;
        ANTENNAMAXAREACAR 41.41  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.42 1.46 8.72 1.74 ;
        RECT  8.34 1.92 8.62 2.52 ;
        RECT  8.34 0.62 8.62 1.22 ;
        RECT  8.42 0.62 8.58 2.52 ;
        END
    END OUT
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.64 1.38 7.94 1.76 ;
        END
    END IN3
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.78 1.42 1.18 1.70 ;
        END
    END IN1
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 8.80 0.28 ;
        RECT  8.34 -0.28 8.62 0.32 ;
        RECT  7.82 0.62 8.10 1.22 ;
        RECT  7.88 -0.28 8.04 1.22 ;
        RECT  1.48 -0.28 1.76 0.58 ;
        RECT  0.72 0.78 1.00 1.06 ;
        RECT  0.78 -0.28 0.94 1.06 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 8.80 3.48 ;
        RECT  8.34 2.88 8.62 3.48 ;
        RECT  7.82 1.92 8.10 2.52 ;
        RECT  7.84 1.92 8.00 3.48 ;
        RECT  1.72 1.92 2.00 2.20 ;
        RECT  1.82 1.92 1.98 3.48 ;
        RECT  0.72 1.86 1.00 2.14 ;
        RECT  0.78 1.86 0.94 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.20 0.78 0.48 1.06 ;
        RECT  0.20 1.86 0.48 2.14 ;
        RECT  0.22 0.78 0.38 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  2.24 0.76 2.52 1.04 ;
        RECT  2.28 1.22 2.66 1.50 ;
        RECT  2.28 0.76 2.44 2.20 ;
        RECT  2.24 1.92 2.52 2.20 ;
        RECT  2.72 0.76 3.00 1.04 ;
        RECT  2.82 0.76 2.98 2.20 ;
        RECT  2.72 1.92 3.00 2.20 ;
        RECT  2.72 1.92 2.88 2.63 ;
        RECT  2.58 2.35 2.88 2.63 ;
        RECT  1.92 0.44 3.92 0.60 ;
        RECT  3.76 0.44 3.92 1.04 ;
        RECT  1.92 0.44 2.08 0.94 ;
        RECT  1.24 0.78 2.08 0.94 ;
        RECT  3.76 0.76 4.04 1.04 ;
        RECT  1.24 0.78 1.52 1.06 ;
        RECT  3.82 0.76 3.98 2.20 ;
        RECT  1.24 1.86 1.52 2.14 ;
        RECT  3.76 1.92 4.04 2.20 ;
        RECT  1.34 0.78 1.50 2.68 ;
        RECT  1.34 2.40 1.66 2.68 ;
        RECT  4.80 0.76 5.08 1.04 ;
        RECT  4.92 1.54 5.22 1.82 ;
        RECT  4.92 0.76 5.08 2.20 ;
        RECT  4.80 1.92 5.08 2.20 ;
        RECT  3.24 0.76 3.52 1.04 ;
        RECT  5.40 0.76 5.68 1.04 ;
        RECT  5.46 0.76 5.62 2.20 ;
        RECT  3.30 0.76 3.46 2.20 ;
        RECT  3.24 1.92 3.52 2.20 ;
        RECT  5.40 1.92 5.68 2.20 ;
        RECT  3.36 1.92 3.52 2.52 ;
        RECT  5.40 1.92 5.56 2.52 ;
        RECT  3.36 2.36 5.56 2.52 ;
        RECT  4.40 0.44 6.60 0.60 ;
        RECT  4.40 0.44 4.56 1.04 ;
        RECT  4.28 0.76 4.56 1.04 ;
        RECT  6.44 0.76 6.72 1.04 ;
        RECT  4.34 0.76 4.50 2.20 ;
        RECT  6.44 0.44 6.60 2.20 ;
        RECT  4.28 1.92 4.56 2.20 ;
        RECT  6.44 1.92 6.72 2.20 ;
        RECT  5.92 0.76 6.20 1.04 ;
        RECT  5.98 0.76 6.14 2.20 ;
        RECT  5.92 1.92 6.20 2.20 ;
        RECT  6.04 1.92 6.20 2.70 ;
        RECT  6.04 2.54 7.42 2.70 ;
        RECT  7.14 2.48 7.42 2.76 ;
        RECT  7.26 0.76 7.54 1.04 ;
        RECT  7.12 1.14 7.42 1.42 ;
        RECT  7.26 0.76 7.42 2.20 ;
        RECT  7.26 1.92 7.54 2.20 ;
    END
END XOR3SP2V1_0

MACRO XOR3SP1V1_0
    CLASS CORE ;
    FOREIGN XOR3SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.78 1.42 1.18 1.70 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.66 1.46 2.10 1.74 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.64 1.34 7.94 1.76 ;
        END
    END IN3
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 16.84  LAYER ME1  ;
        ANTENNADIFFAREA 6.45  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.34  LAYER ME1  ;
        ANTENNAMAXAREACAR 50.12  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.42 1.46 8.72 1.74 ;
        RECT  8.30 1.92 8.58 2.20 ;
        RECT  8.42 0.76 8.58 2.20 ;
        RECT  8.30 0.76 8.58 1.04 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 8.80 3.48 ;
        RECT  8.34 2.88 8.62 3.48 ;
        RECT  7.78 1.92 8.06 2.20 ;
        RECT  7.84 1.92 8.00 3.48 ;
        RECT  1.72 1.92 2.00 2.20 ;
        RECT  1.82 1.92 1.98 3.48 ;
        RECT  0.72 1.86 1.00 2.14 ;
        RECT  0.78 1.86 0.94 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 8.80 0.28 ;
        RECT  8.34 -0.28 8.62 0.32 ;
        RECT  7.78 0.76 8.06 1.04 ;
        RECT  7.84 -0.28 8.00 1.04 ;
        RECT  1.48 -0.28 1.76 0.58 ;
        RECT  0.72 0.78 1.00 1.06 ;
        RECT  0.78 -0.28 0.94 1.06 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.20 0.78 0.48 1.06 ;
        RECT  0.20 1.86 0.48 2.14 ;
        RECT  0.22 0.78 0.38 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  2.24 0.76 2.52 1.04 ;
        RECT  2.28 1.22 2.66 1.50 ;
        RECT  2.28 0.76 2.44 2.20 ;
        RECT  2.24 1.92 2.52 2.20 ;
        RECT  2.72 0.76 3.00 1.04 ;
        RECT  2.82 0.76 2.98 2.20 ;
        RECT  2.72 1.92 3.00 2.20 ;
        RECT  2.72 1.92 2.88 2.63 ;
        RECT  2.58 2.35 2.88 2.63 ;
        RECT  1.92 0.44 3.92 0.60 ;
        RECT  3.76 0.44 3.92 1.04 ;
        RECT  1.92 0.44 2.08 0.94 ;
        RECT  1.24 0.78 2.08 0.94 ;
        RECT  3.76 0.76 4.04 1.04 ;
        RECT  1.24 0.78 1.52 1.06 ;
        RECT  3.82 0.76 3.98 2.20 ;
        RECT  1.24 1.86 1.52 2.14 ;
        RECT  3.76 1.92 4.04 2.20 ;
        RECT  1.34 0.78 1.50 2.68 ;
        RECT  1.34 2.40 1.66 2.68 ;
        RECT  4.80 0.76 5.08 1.04 ;
        RECT  4.92 1.54 5.22 1.82 ;
        RECT  4.92 0.76 5.08 2.20 ;
        RECT  4.80 1.92 5.08 2.20 ;
        RECT  3.24 0.76 3.52 1.04 ;
        RECT  5.40 0.76 5.68 1.04 ;
        RECT  5.46 0.76 5.62 2.20 ;
        RECT  3.30 0.76 3.46 2.20 ;
        RECT  3.24 1.92 3.52 2.20 ;
        RECT  5.40 1.92 5.68 2.20 ;
        RECT  3.36 1.92 3.52 2.52 ;
        RECT  5.40 1.92 5.56 2.52 ;
        RECT  3.36 2.36 5.56 2.52 ;
        RECT  4.40 0.44 6.60 0.60 ;
        RECT  4.40 0.44 4.56 1.04 ;
        RECT  4.28 0.76 4.56 1.04 ;
        RECT  6.44 0.76 6.72 1.04 ;
        RECT  4.34 0.76 4.50 2.20 ;
        RECT  6.44 0.44 6.60 2.20 ;
        RECT  4.28 1.92 4.56 2.20 ;
        RECT  6.44 1.92 6.72 2.20 ;
        RECT  5.92 0.76 6.20 1.04 ;
        RECT  5.98 0.76 6.14 2.20 ;
        RECT  5.92 1.92 6.20 2.20 ;
        RECT  6.04 1.92 6.20 2.70 ;
        RECT  6.04 2.54 7.42 2.70 ;
        RECT  7.14 2.48 7.42 2.76 ;
        RECT  7.26 0.76 7.54 1.04 ;
        RECT  7.12 1.14 7.42 1.42 ;
        RECT  7.26 0.76 7.42 2.20 ;
        RECT  7.26 1.92 7.54 2.20 ;
    END
END XOR3SP1V1_0

MACRO XOR2SP8V1_0
    CLASS CORE ;
    FOREIGN XOR2SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.90 1.26 1.18 1.68 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.42 1.12 0.70 1.54 ;
        END
    END IN2
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 10.90  LAYER ME1  ;
        ANTENNADIFFAREA 5.85  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.71  LAYER ME1  ;
        ANTENNAMAXAREACAR 15.35  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.06 1.84 5.34 2.12 ;
        RECT  5.06 0.96 5.34 1.24 ;
        RECT  5.06 0.96 5.22 2.12 ;
        RECT  4.12 1.52 5.22 1.68 ;
        RECT  4.02 1.84 4.30 2.12 ;
        RECT  4.02 0.96 4.30 1.24 ;
        RECT  4.12 0.96 4.28 2.12 ;
        END
    END OUT
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 6.00 0.28 ;
        RECT  5.58 0.64 5.86 0.92 ;
        RECT  5.54 -0.28 5.82 0.32 ;
        RECT  5.64 -0.28 5.80 0.92 ;
        RECT  4.54 0.64 4.82 0.92 ;
        RECT  4.60 -0.28 4.76 0.92 ;
        RECT  3.50 0.64 3.78 0.92 ;
        RECT  3.52 -0.28 3.68 0.92 ;
        RECT  0.76 0.68 1.04 0.96 ;
        RECT  0.82 -0.28 0.98 0.96 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 6.00 3.48 ;
        RECT  5.58 2.16 5.86 2.44 ;
        RECT  5.54 2.88 5.82 3.48 ;
        RECT  5.64 2.16 5.80 3.48 ;
        RECT  4.54 2.16 4.82 2.44 ;
        RECT  4.60 2.16 4.76 3.48 ;
        RECT  3.50 2.16 3.78 2.44 ;
        RECT  3.56 2.16 3.72 3.48 ;
        RECT  0.76 1.84 1.04 2.12 ;
        RECT  0.82 1.84 0.98 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.68 0.52 0.96 ;
        RECT  0.10 1.84 0.52 2.12 ;
        RECT  0.10 0.68 0.26 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  1.92 0.44 3.08 0.60 ;
        RECT  2.80 0.44 3.08 0.72 ;
        RECT  1.92 0.44 2.08 0.96 ;
        RECT  1.80 0.68 2.08 0.96 ;
        RECT  1.86 0.68 2.02 2.12 ;
        RECT  1.80 1.84 2.08 2.12 ;
        RECT  2.36 0.76 2.64 1.04 ;
        RECT  2.94 0.96 3.22 1.24 ;
        RECT  2.38 1.46 3.16 1.62 ;
        RECT  2.38 0.76 2.54 2.12 ;
        RECT  3.00 0.96 3.16 2.12 ;
        RECT  2.32 1.84 2.60 2.12 ;
        RECT  2.94 1.84 3.22 2.12 ;
        RECT  1.28 0.68 1.56 0.96 ;
        RECT  1.34 0.68 1.50 2.12 ;
        RECT  1.28 1.84 1.56 2.12 ;
        RECT  1.40 1.84 1.56 2.44 ;
        RECT  1.40 2.28 3.34 2.44 ;
        RECT  3.06 2.28 3.34 2.56 ;
    END
END XOR2SP8V1_0

MACRO XOR2SP4V1_0
    CLASS CORE ;
    FOREIGN XOR2SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 9.10  LAYER ME1  ;
        ANTENNADIFFAREA 4.43  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.42  LAYER ME1  ;
        ANTENNAMAXAREACAR 21.53  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.02 1.84 4.30 2.12 ;
        RECT  4.02 0.96 4.30 1.24 ;
        RECT  4.12 0.96 4.28 2.12 ;
        END
    END OUT
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.42 1.12 0.70 1.54 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.90 1.26 1.18 1.68 ;
        END
    END IN1
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 5.20 0.28 ;
        RECT  4.60 -0.28 5.02 0.32 ;
        RECT  4.54 0.64 4.82 0.92 ;
        RECT  4.60 -0.28 4.76 0.92 ;
        RECT  3.50 0.64 3.78 0.92 ;
        RECT  3.52 -0.28 3.68 0.92 ;
        RECT  0.76 0.68 1.04 0.96 ;
        RECT  0.82 -0.28 0.98 0.96 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 5.20 3.48 ;
        RECT  4.60 2.88 5.02 3.48 ;
        RECT  4.54 2.16 4.82 2.44 ;
        RECT  4.60 2.16 4.76 3.48 ;
        RECT  3.50 2.16 3.78 2.44 ;
        RECT  3.56 2.16 3.72 3.48 ;
        RECT  0.76 1.84 1.04 2.12 ;
        RECT  0.82 1.84 0.98 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.68 0.52 0.96 ;
        RECT  0.10 1.84 0.52 2.12 ;
        RECT  0.10 0.68 0.26 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  1.92 0.44 3.08 0.60 ;
        RECT  2.80 0.44 3.08 0.72 ;
        RECT  1.92 0.44 2.08 0.96 ;
        RECT  1.80 0.68 2.08 0.96 ;
        RECT  1.86 0.68 2.02 2.12 ;
        RECT  1.80 1.84 2.08 2.12 ;
        RECT  2.36 0.76 2.64 1.04 ;
        RECT  2.94 0.96 3.22 1.24 ;
        RECT  2.38 1.46 3.16 1.62 ;
        RECT  2.38 0.76 2.54 2.12 ;
        RECT  3.00 0.96 3.16 2.12 ;
        RECT  2.32 1.84 2.60 2.12 ;
        RECT  2.94 1.84 3.22 2.12 ;
        RECT  1.28 0.68 1.56 0.96 ;
        RECT  1.34 0.68 1.50 2.12 ;
        RECT  1.28 1.84 1.56 2.12 ;
        RECT  1.40 1.84 1.56 2.44 ;
        RECT  1.40 2.28 3.34 2.44 ;
        RECT  3.06 2.28 3.34 2.56 ;
    END
END XOR2SP4V1_0

MACRO XOR2SP2V1_0
    CLASS CORE ;
    FOREIGN XOR2SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 7.91  LAYER ME1  ;
        ANTENNADIFFAREA 3.69  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.28  LAYER ME1  ;
        ANTENNAMAXAREACAR 28.41  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.02 1.84 4.30 2.12 ;
        RECT  4.02 0.96 4.30 1.24 ;
        RECT  4.12 0.96 4.28 2.12 ;
        END
    END OUT
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.90 1.26 1.18 1.68 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.42 1.12 0.70 1.54 ;
        END
    END IN2
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.40 0.28 ;
        RECT  3.94 -0.28 4.22 0.32 ;
        RECT  3.50 0.64 3.78 0.92 ;
        RECT  3.52 -0.28 3.68 0.92 ;
        RECT  0.76 0.68 1.04 0.96 ;
        RECT  0.82 -0.28 0.98 0.96 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.40 3.48 ;
        RECT  3.94 2.88 4.22 3.48 ;
        RECT  3.50 2.16 3.78 2.44 ;
        RECT  3.56 2.16 3.72 3.48 ;
        RECT  0.76 1.84 1.04 2.12 ;
        RECT  0.82 1.84 0.98 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.68 0.52 0.96 ;
        RECT  0.10 1.84 0.52 2.12 ;
        RECT  0.10 0.68 0.26 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  1.92 0.44 3.08 0.60 ;
        RECT  2.80 0.44 3.08 0.72 ;
        RECT  1.92 0.44 2.08 0.96 ;
        RECT  1.80 0.68 2.08 0.96 ;
        RECT  1.86 0.68 2.02 2.12 ;
        RECT  1.80 1.84 2.08 2.12 ;
        RECT  2.36 0.76 2.64 1.04 ;
        RECT  2.94 0.96 3.22 1.24 ;
        RECT  2.38 1.46 3.16 1.62 ;
        RECT  2.38 0.76 2.54 2.12 ;
        RECT  3.00 0.96 3.16 2.12 ;
        RECT  2.32 1.84 2.60 2.12 ;
        RECT  2.94 1.84 3.22 2.12 ;
        RECT  1.28 0.68 1.56 0.96 ;
        RECT  1.34 0.68 1.50 2.12 ;
        RECT  1.28 1.84 1.56 2.12 ;
        RECT  1.40 1.84 1.56 2.44 ;
        RECT  1.40 2.28 3.34 2.44 ;
        RECT  3.06 2.28 3.34 2.56 ;
    END
END XOR2SP2V1_0

MACRO XOR2SP1V1_0
    CLASS CORE ;
    FOREIGN XOR2SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.90 1.26 1.18 1.68 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.42 1.12 0.70 1.54 ;
        END
    END IN2
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 8.02  LAYER ME1  ;
        ANTENNADIFFAREA 3.23  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        ANTENNAMAXAREACAR 39.79  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.98 1.84 4.28 2.12 ;
        RECT  4.12 0.96 4.28 2.12 ;
        RECT  3.98 0.96 4.28 1.24 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.40 3.48 ;
        RECT  3.94 2.88 4.22 3.48 ;
        RECT  3.46 1.84 3.74 2.12 ;
        RECT  3.56 1.84 3.72 3.48 ;
        RECT  0.76 1.84 1.04 2.12 ;
        RECT  0.82 1.84 0.98 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.40 0.28 ;
        RECT  3.94 -0.28 4.22 0.32 ;
        RECT  3.46 0.96 3.74 1.24 ;
        RECT  3.52 -0.28 3.68 1.24 ;
        RECT  0.76 0.68 1.04 0.96 ;
        RECT  0.82 -0.28 0.98 0.96 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.68 0.52 0.96 ;
        RECT  0.10 1.84 0.52 2.12 ;
        RECT  0.10 0.68 0.26 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  1.92 0.44 3.08 0.60 ;
        RECT  2.80 0.44 3.08 0.72 ;
        RECT  1.92 0.44 2.08 0.96 ;
        RECT  1.80 0.68 2.08 0.96 ;
        RECT  1.86 0.68 2.02 2.12 ;
        RECT  1.80 1.84 2.08 2.12 ;
        RECT  2.36 0.76 2.64 1.04 ;
        RECT  2.94 0.96 3.22 1.24 ;
        RECT  2.38 1.46 3.16 1.62 ;
        RECT  2.38 0.76 2.54 2.12 ;
        RECT  3.00 0.96 3.16 2.12 ;
        RECT  2.32 1.84 2.60 2.12 ;
        RECT  2.94 1.84 3.22 2.12 ;
        RECT  1.28 0.68 1.56 0.96 ;
        RECT  1.34 0.68 1.50 2.12 ;
        RECT  1.28 1.84 1.56 2.12 ;
        RECT  1.40 1.84 1.56 2.44 ;
        RECT  1.40 2.28 3.40 2.44 ;
        RECT  3.12 2.28 3.40 2.56 ;
    END
END XOR2SP1V1_0

MACRO XNR3SP8V1_0
    CLASS CORE ;
    FOREIGN XNR3SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 20.39  LAYER ME1  ;
        ANTENNADIFFAREA 9.43  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.84  LAYER ME1  ;
        ANTENNAMAXAREACAR 24.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.44 1.92 9.72 2.52 ;
        RECT  9.44 0.64 9.72 1.24 ;
        RECT  9.44 0.64 9.60 2.52 ;
        RECT  8.46 1.52 9.60 1.68 ;
        RECT  8.46 1.46 8.74 1.74 ;
        RECT  8.40 1.92 8.68 2.52 ;
        RECT  8.46 0.64 8.68 2.52 ;
        RECT  8.40 0.64 8.68 1.24 ;
        END
    END OUT
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.66 1.44 8.05 1.76 ;
        END
    END IN3
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.78 1.42 1.18 1.70 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.66 1.46 2.10 1.74 ;
        END
    END IN2
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 10.40 0.28 ;
        RECT  9.96 0.64 10.24 1.24 ;
        RECT  9.94 -0.28 10.22 0.32 ;
        RECT  10.02 -0.28 10.18 1.24 ;
        RECT  8.92 0.64 9.20 1.24 ;
        RECT  8.98 -0.28 9.14 1.24 ;
        RECT  7.88 0.64 8.16 1.24 ;
        RECT  7.94 -0.28 8.10 1.24 ;
        RECT  1.72 0.76 2.00 1.04 ;
        RECT  1.78 -0.28 1.94 1.04 ;
        RECT  0.72 0.78 1.00 1.06 ;
        RECT  0.78 -0.28 0.94 1.06 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 10.40 3.48 ;
        RECT  9.96 1.92 10.24 2.52 ;
        RECT  9.94 2.88 10.22 3.48 ;
        RECT  10.02 1.92 10.18 3.48 ;
        RECT  8.92 1.92 9.20 2.52 ;
        RECT  8.98 1.92 9.14 3.48 ;
        RECT  7.88 1.92 8.16 2.52 ;
        RECT  7.94 1.92 8.10 3.48 ;
        RECT  1.72 1.92 2.00 2.20 ;
        RECT  1.82 1.92 1.98 3.48 ;
        RECT  0.72 1.86 1.00 2.14 ;
        RECT  0.78 1.86 0.94 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.20 0.78 0.48 1.06 ;
        RECT  0.20 1.86 0.48 2.14 ;
        RECT  0.22 0.78 0.38 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  1.24 0.78 1.52 1.06 ;
        RECT  1.24 1.86 1.52 2.14 ;
        RECT  1.34 0.78 1.50 2.70 ;
        RECT  1.34 2.42 1.66 2.70 ;
        RECT  2.24 0.76 2.52 1.04 ;
        RECT  2.36 1.12 2.94 1.40 ;
        RECT  2.36 0.76 2.52 2.20 ;
        RECT  2.24 1.92 2.52 2.20 ;
        RECT  3.12 0.76 3.40 1.04 ;
        RECT  3.22 0.76 3.38 2.20 ;
        RECT  2.68 1.92 3.40 2.20 ;
        RECT  4.16 0.76 4.44 1.04 ;
        RECT  4.22 0.76 4.38 2.20 ;
        RECT  4.16 1.92 4.44 2.20 ;
        RECT  4.16 1.92 4.32 2.68 ;
        RECT  2.38 2.52 4.32 2.68 ;
        RECT  2.38 2.42 2.66 2.70 ;
        RECT  5.20 0.76 5.48 1.04 ;
        RECT  5.32 1.54 5.62 1.82 ;
        RECT  5.32 0.76 5.48 2.20 ;
        RECT  5.20 1.92 5.48 2.20 ;
        RECT  4.68 0.76 4.96 1.04 ;
        RECT  5.80 0.76 6.08 1.04 ;
        RECT  5.86 0.76 6.02 2.20 ;
        RECT  4.74 0.76 4.90 2.20 ;
        RECT  4.68 1.92 4.96 2.20 ;
        RECT  5.80 1.92 6.08 2.20 ;
        RECT  4.80 1.92 4.96 2.52 ;
        RECT  5.80 1.92 5.96 2.52 ;
        RECT  4.80 2.36 5.96 2.52 ;
        RECT  3.76 0.44 7.00 0.60 ;
        RECT  3.76 0.44 3.92 1.04 ;
        RECT  3.64 0.76 3.92 1.04 ;
        RECT  6.84 0.76 7.12 1.04 ;
        RECT  3.70 0.76 3.86 2.20 ;
        RECT  6.84 0.44 7.00 2.20 ;
        RECT  3.64 1.92 3.92 2.20 ;
        RECT  6.84 1.92 7.12 2.20 ;
        RECT  6.32 0.76 6.60 1.04 ;
        RECT  6.38 0.76 6.54 2.20 ;
        RECT  6.32 1.92 6.60 2.20 ;
        RECT  6.44 1.92 6.60 2.70 ;
        RECT  6.44 2.54 7.48 2.70 ;
        RECT  7.20 2.48 7.48 2.76 ;
        RECT  7.32 0.76 7.60 1.04 ;
        RECT  7.18 1.19 7.48 1.47 ;
        RECT  7.32 0.76 7.48 2.20 ;
        RECT  7.32 1.92 7.60 2.20 ;
    END
END XNR3SP8V1_0

MACRO XNR3SP4V1_0
    CLASS CORE ;
    FOREIGN XNR3SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.66 1.46 2.10 1.74 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.78 1.42 1.18 1.70 ;
        END
    END IN1
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.66 1.44 8.05 1.76 ;
        END
    END IN3
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 18.48  LAYER ME1  ;
        ANTENNADIFFAREA 7.74  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.56  LAYER ME1  ;
        ANTENNAMAXAREACAR 33.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.46 1.46 8.72 1.74 ;
        RECT  8.40 1.92 8.68 2.52 ;
        RECT  8.46 0.64 8.68 2.52 ;
        RECT  8.40 0.64 8.68 1.24 ;
        END
    END OUT
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 9.60 0.28 ;
        RECT  8.98 -0.28 9.42 0.32 ;
        RECT  8.92 0.64 9.20 1.24 ;
        RECT  8.98 -0.28 9.14 1.24 ;
        RECT  7.88 0.64 8.16 1.24 ;
        RECT  7.94 -0.28 8.10 1.24 ;
        RECT  1.72 0.76 2.00 1.04 ;
        RECT  1.78 -0.28 1.94 1.04 ;
        RECT  0.72 0.78 1.00 1.06 ;
        RECT  0.78 -0.28 0.94 1.06 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 9.60 3.48 ;
        RECT  8.98 2.88 9.42 3.48 ;
        RECT  8.92 1.92 9.20 2.52 ;
        RECT  8.98 1.92 9.14 3.48 ;
        RECT  7.88 1.92 8.16 2.52 ;
        RECT  7.94 1.92 8.10 3.48 ;
        RECT  1.72 1.92 2.00 2.20 ;
        RECT  1.82 1.92 1.98 3.48 ;
        RECT  0.72 1.86 1.00 2.14 ;
        RECT  0.78 1.86 0.94 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.20 0.78 0.48 1.06 ;
        RECT  0.20 1.86 0.48 2.14 ;
        RECT  0.22 0.78 0.38 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  1.24 0.78 1.52 1.06 ;
        RECT  1.24 1.86 1.52 2.14 ;
        RECT  1.34 0.78 1.50 2.68 ;
        RECT  1.38 2.42 1.66 2.70 ;
        RECT  2.24 0.76 2.52 1.04 ;
        RECT  2.36 1.12 2.94 1.40 ;
        RECT  2.36 0.76 2.52 2.20 ;
        RECT  2.24 1.92 2.52 2.20 ;
        RECT  3.12 0.76 3.40 1.04 ;
        RECT  3.22 0.76 3.38 2.20 ;
        RECT  2.68 1.92 3.40 2.20 ;
        RECT  4.16 0.76 4.44 1.04 ;
        RECT  4.22 0.76 4.38 2.20 ;
        RECT  4.16 1.92 4.44 2.20 ;
        RECT  4.16 1.92 4.32 2.68 ;
        RECT  2.38 2.52 4.32 2.68 ;
        RECT  2.38 2.42 2.66 2.70 ;
        RECT  5.20 0.76 5.48 1.04 ;
        RECT  5.32 1.54 5.62 1.82 ;
        RECT  5.32 0.76 5.48 2.20 ;
        RECT  5.20 1.92 5.48 2.20 ;
        RECT  4.68 0.76 4.96 1.04 ;
        RECT  5.80 0.76 6.08 1.04 ;
        RECT  5.86 0.76 6.02 2.20 ;
        RECT  4.74 0.76 4.90 2.20 ;
        RECT  4.68 1.92 4.96 2.20 ;
        RECT  5.80 1.92 6.08 2.20 ;
        RECT  4.80 1.92 4.96 2.52 ;
        RECT  5.80 1.92 5.96 2.52 ;
        RECT  4.80 2.36 5.96 2.52 ;
        RECT  3.76 0.44 7.00 0.60 ;
        RECT  3.76 0.44 3.92 1.04 ;
        RECT  3.64 0.76 3.92 1.04 ;
        RECT  6.84 0.76 7.12 1.04 ;
        RECT  3.70 0.76 3.86 2.20 ;
        RECT  6.84 0.44 7.00 2.20 ;
        RECT  3.64 1.92 3.92 2.20 ;
        RECT  6.84 1.92 7.12 2.20 ;
        RECT  6.32 0.76 6.60 1.04 ;
        RECT  6.38 0.76 6.54 2.20 ;
        RECT  6.32 1.92 6.60 2.20 ;
        RECT  6.44 1.92 6.60 2.70 ;
        RECT  6.44 2.54 7.48 2.70 ;
        RECT  7.20 2.48 7.48 2.76 ;
        RECT  7.32 0.76 7.60 1.04 ;
        RECT  7.18 1.19 7.48 1.47 ;
        RECT  7.32 0.76 7.48 2.20 ;
        RECT  7.32 1.92 7.60 2.20 ;
    END
END XNR3SP4V1_0

MACRO XNR3SP2V1_0
    CLASS CORE ;
    FOREIGN XNR3SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 17.13  LAYER ME1  ;
        ANTENNADIFFAREA 6.77  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.41  LAYER ME1  ;
        ANTENNAMAXAREACAR 41.50  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.46 1.46 8.72 1.74 ;
        RECT  8.40 1.92 8.68 2.52 ;
        RECT  8.46 0.64 8.68 2.52 ;
        RECT  8.40 0.64 8.68 1.24 ;
        END
    END OUT
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.66 1.44 8.05 1.76 ;
        END
    END IN3
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.78 1.42 1.18 1.70 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.66 1.46 2.10 1.74 ;
        END
    END IN2
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 8.80 3.48 ;
        RECT  8.34 2.88 8.62 3.48 ;
        RECT  7.88 1.92 8.16 2.52 ;
        RECT  7.94 1.92 8.10 3.48 ;
        RECT  1.72 1.92 2.00 2.20 ;
        RECT  1.82 1.92 1.98 3.48 ;
        RECT  0.72 1.86 1.00 2.14 ;
        RECT  0.78 1.86 0.94 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 8.80 0.28 ;
        RECT  8.34 -0.28 8.62 0.32 ;
        RECT  7.88 0.64 8.16 1.24 ;
        RECT  7.94 -0.28 8.10 1.24 ;
        RECT  1.72 0.76 2.00 1.04 ;
        RECT  1.78 -0.28 1.94 1.04 ;
        RECT  0.72 0.78 1.00 1.06 ;
        RECT  0.78 -0.28 0.94 1.06 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.20 0.78 0.48 1.06 ;
        RECT  0.20 1.86 0.48 2.14 ;
        RECT  0.22 0.78 0.38 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  1.24 0.78 1.52 1.06 ;
        RECT  1.24 1.86 1.52 2.14 ;
        RECT  1.34 0.78 1.50 2.70 ;
        RECT  1.34 2.42 1.66 2.70 ;
        RECT  2.24 0.76 2.52 1.04 ;
        RECT  2.36 1.12 2.94 1.40 ;
        RECT  2.36 0.76 2.52 2.20 ;
        RECT  2.24 1.92 2.52 2.20 ;
        RECT  3.12 0.76 3.40 1.04 ;
        RECT  3.22 0.76 3.38 2.20 ;
        RECT  2.68 1.92 3.40 2.20 ;
        RECT  4.16 0.76 4.44 1.04 ;
        RECT  4.22 0.76 4.38 2.20 ;
        RECT  4.16 1.92 4.44 2.20 ;
        RECT  4.16 1.92 4.32 2.68 ;
        RECT  2.38 2.52 4.32 2.68 ;
        RECT  2.38 2.42 2.66 2.70 ;
        RECT  5.20 0.76 5.48 1.04 ;
        RECT  5.32 1.54 5.62 1.82 ;
        RECT  5.32 0.76 5.48 2.20 ;
        RECT  5.20 1.92 5.48 2.20 ;
        RECT  4.68 0.76 4.96 1.04 ;
        RECT  5.80 0.76 6.08 1.04 ;
        RECT  5.86 0.76 6.02 2.20 ;
        RECT  4.74 0.76 4.90 2.20 ;
        RECT  4.68 1.92 4.96 2.20 ;
        RECT  5.80 1.92 6.08 2.20 ;
        RECT  4.80 1.92 4.96 2.52 ;
        RECT  5.80 1.92 5.96 2.52 ;
        RECT  4.80 2.36 5.96 2.52 ;
        RECT  3.76 0.44 7.00 0.60 ;
        RECT  3.76 0.44 3.92 1.04 ;
        RECT  3.64 0.76 3.92 1.04 ;
        RECT  6.84 0.76 7.12 1.04 ;
        RECT  3.70 0.76 3.86 2.20 ;
        RECT  6.84 0.44 7.00 2.20 ;
        RECT  3.64 1.92 3.92 2.20 ;
        RECT  6.84 1.92 7.12 2.20 ;
        RECT  6.32 0.76 6.60 1.04 ;
        RECT  6.38 0.76 6.54 2.20 ;
        RECT  6.32 1.92 6.60 2.20 ;
        RECT  6.44 1.92 6.60 2.70 ;
        RECT  6.44 2.54 7.48 2.70 ;
        RECT  7.20 2.48 7.48 2.76 ;
        RECT  7.32 0.76 7.60 1.04 ;
        RECT  7.18 1.19 7.48 1.47 ;
        RECT  7.32 0.76 7.48 2.20 ;
        RECT  7.32 1.92 7.60 2.20 ;
    END
END XNR3SP2V1_0

MACRO XNR3SP1V1_0
    CLASS CORE ;
    FOREIGN XNR3SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.66 1.46 2.10 1.74 ;
        END
    END IN2
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 16.86  LAYER ME1  ;
        ANTENNADIFFAREA 6.31  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.34  LAYER ME1  ;
        ANTENNAMAXAREACAR 50.19  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.46 1.46 8.72 1.74 ;
        RECT  8.36 1.92 8.64 2.20 ;
        RECT  8.46 0.76 8.64 2.20 ;
        RECT  8.36 0.76 8.64 1.04 ;
        END
    END OUT
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.66 1.34 7.96 1.76 ;
        END
    END IN3
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.78 1.42 1.18 1.70 ;
        END
    END IN1
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 8.80 3.48 ;
        RECT  8.34 2.88 8.62 3.48 ;
        RECT  7.84 1.92 8.12 2.20 ;
        RECT  7.90 1.92 8.06 3.48 ;
        RECT  1.72 1.92 2.00 2.20 ;
        RECT  1.82 1.92 1.98 3.48 ;
        RECT  0.72 1.86 1.00 2.14 ;
        RECT  0.78 1.86 0.94 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 8.80 0.28 ;
        RECT  8.34 -0.28 8.62 0.32 ;
        RECT  7.84 0.76 8.12 1.04 ;
        RECT  7.90 -0.28 8.06 1.04 ;
        RECT  1.72 0.76 2.00 1.04 ;
        RECT  1.78 -0.28 1.94 1.04 ;
        RECT  0.72 0.78 1.00 1.06 ;
        RECT  0.78 -0.28 0.94 1.06 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.20 0.78 0.48 1.06 ;
        RECT  0.20 1.86 0.48 2.14 ;
        RECT  0.22 0.78 0.38 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  1.24 0.78 1.52 1.06 ;
        RECT  1.24 1.86 1.52 2.14 ;
        RECT  1.34 0.78 1.50 2.70 ;
        RECT  1.34 2.42 1.66 2.70 ;
        RECT  2.24 0.76 2.52 1.04 ;
        RECT  2.36 1.12 2.94 1.40 ;
        RECT  2.36 0.76 2.52 2.20 ;
        RECT  2.24 1.92 2.52 2.20 ;
        RECT  3.12 0.76 3.40 1.04 ;
        RECT  3.22 0.76 3.38 2.20 ;
        RECT  2.68 1.92 3.40 2.20 ;
        RECT  4.16 0.76 4.44 1.04 ;
        RECT  4.22 0.76 4.38 2.20 ;
        RECT  4.16 1.92 4.44 2.20 ;
        RECT  4.16 1.92 4.32 2.68 ;
        RECT  2.38 2.52 4.32 2.68 ;
        RECT  2.38 2.42 2.66 2.70 ;
        RECT  5.20 0.76 5.48 1.04 ;
        RECT  5.32 1.54 5.62 1.82 ;
        RECT  5.32 0.76 5.48 2.20 ;
        RECT  5.20 1.92 5.48 2.20 ;
        RECT  4.68 0.76 4.96 1.04 ;
        RECT  5.80 0.76 6.08 1.04 ;
        RECT  5.86 0.76 6.02 2.20 ;
        RECT  4.74 0.76 4.90 2.20 ;
        RECT  4.68 1.92 4.96 2.20 ;
        RECT  5.80 1.92 6.08 2.20 ;
        RECT  4.80 1.92 4.96 2.52 ;
        RECT  5.80 1.92 5.96 2.52 ;
        RECT  4.80 2.36 5.96 2.52 ;
        RECT  3.76 0.44 7.00 0.60 ;
        RECT  3.76 0.44 3.92 1.04 ;
        RECT  3.64 0.76 3.92 1.04 ;
        RECT  6.84 0.76 7.12 1.04 ;
        RECT  3.70 0.76 3.86 2.20 ;
        RECT  6.84 0.44 7.00 2.20 ;
        RECT  3.64 1.92 3.92 2.20 ;
        RECT  6.84 1.92 7.12 2.20 ;
        RECT  6.32 0.76 6.60 1.04 ;
        RECT  6.38 0.76 6.54 2.20 ;
        RECT  6.32 1.92 6.60 2.20 ;
        RECT  6.44 1.92 6.60 2.70 ;
        RECT  6.44 2.54 7.48 2.70 ;
        RECT  7.20 2.48 7.48 2.76 ;
        RECT  7.32 0.76 7.60 1.04 ;
        RECT  7.18 1.19 7.48 1.47 ;
        RECT  7.32 0.76 7.48 2.20 ;
        RECT  7.32 1.92 7.60 2.20 ;
    END
END XNR3SP1V1_0

MACRO XNR2SP8V1_0
    CLASS CORE ;
    FOREIGN XNR2SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 10.99  LAYER ME1  ;
        ANTENNADIFFAREA 5.88  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.74  LAYER ME1  ;
        ANTENNAMAXAREACAR 14.77  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.06 1.84 5.34 2.12 ;
        RECT  5.06 0.96 5.34 1.24 ;
        RECT  5.06 0.96 5.22 2.12 ;
        RECT  4.12 1.52 5.22 1.68 ;
        RECT  4.02 1.84 4.30 2.12 ;
        RECT  4.02 0.96 4.30 1.24 ;
        RECT  4.12 0.96 4.28 2.12 ;
        END
    END OUT
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.90 1.33 1.18 1.75 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.42 1.12 0.74 1.54 ;
        END
    END IN2
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 6.00 0.28 ;
        RECT  5.58 0.64 5.86 0.92 ;
        RECT  5.54 -0.28 5.82 0.32 ;
        RECT  5.64 -0.28 5.80 0.92 ;
        RECT  4.54 0.64 4.82 0.92 ;
        RECT  4.60 -0.28 4.76 0.92 ;
        RECT  3.50 0.64 3.78 0.92 ;
        RECT  3.56 -0.28 3.72 0.92 ;
        RECT  0.76 0.68 1.04 0.96 ;
        RECT  0.82 -0.28 0.98 0.96 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 6.00 3.48 ;
        RECT  5.58 2.16 5.86 2.44 ;
        RECT  5.54 2.88 5.82 3.48 ;
        RECT  5.64 2.16 5.80 3.48 ;
        RECT  4.54 2.16 4.82 2.44 ;
        RECT  4.60 2.16 4.76 3.48 ;
        RECT  3.50 1.84 3.78 2.12 ;
        RECT  3.56 1.84 3.72 3.48 ;
        RECT  0.76 1.96 1.04 2.24 ;
        RECT  0.82 1.96 0.98 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.68 0.52 0.96 ;
        RECT  0.10 1.96 0.52 2.24 ;
        RECT  0.10 0.68 0.26 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  1.92 0.44 3.08 0.60 ;
        RECT  2.80 0.44 3.08 0.72 ;
        RECT  1.92 0.44 2.08 0.96 ;
        RECT  1.80 0.68 2.08 0.96 ;
        RECT  1.86 0.68 2.02 2.24 ;
        RECT  1.80 1.96 2.08 2.24 ;
        RECT  2.36 0.76 2.64 1.04 ;
        RECT  2.94 0.96 3.22 1.24 ;
        RECT  2.40 1.46 3.10 1.62 ;
        RECT  2.94 0.96 3.10 2.12 ;
        RECT  2.40 0.76 2.56 2.24 ;
        RECT  2.94 1.84 3.22 2.12 ;
        RECT  2.32 1.96 2.60 2.24 ;
        RECT  1.28 0.68 1.56 0.96 ;
        RECT  1.34 0.68 1.50 2.24 ;
        RECT  1.28 1.96 1.56 2.24 ;
        RECT  1.40 1.96 1.56 2.56 ;
        RECT  3.12 2.28 3.40 2.56 ;
        RECT  1.40 2.40 3.40 2.56 ;
    END
END XNR2SP8V1_0

MACRO XNR2SP4V1_0
    CLASS CORE ;
    FOREIGN XNR2SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.42 1.12 0.74 1.54 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.90 1.33 1.18 1.75 ;
        END
    END IN1
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 9.18  LAYER ME1  ;
        ANTENNADIFFAREA 4.43  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.46  LAYER ME1  ;
        ANTENNAMAXAREACAR 20.14  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.02 1.84 4.30 2.12 ;
        RECT  4.02 0.96 4.30 1.24 ;
        RECT  4.12 0.96 4.28 2.12 ;
        END
    END OUT
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 5.20 0.28 ;
        RECT  4.60 -0.28 5.02 0.32 ;
        RECT  4.54 0.64 4.82 0.92 ;
        RECT  4.60 -0.28 4.76 0.92 ;
        RECT  3.50 0.64 3.78 0.92 ;
        RECT  3.56 -0.28 3.72 0.92 ;
        RECT  0.76 0.68 1.04 0.96 ;
        RECT  0.82 -0.28 0.98 0.96 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 5.20 3.48 ;
        RECT  4.60 2.88 5.02 3.48 ;
        RECT  4.54 2.16 4.82 2.44 ;
        RECT  4.60 2.16 4.76 3.48 ;
        RECT  3.50 1.84 3.78 2.12 ;
        RECT  3.56 1.84 3.72 3.48 ;
        RECT  0.76 1.96 1.04 2.24 ;
        RECT  0.82 1.96 0.98 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.68 0.52 0.96 ;
        RECT  0.10 1.96 0.52 2.24 ;
        RECT  0.10 0.68 0.26 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  1.92 0.44 3.08 0.60 ;
        RECT  2.80 0.44 3.08 0.72 ;
        RECT  1.92 0.44 2.08 0.96 ;
        RECT  1.80 0.68 2.08 0.96 ;
        RECT  1.86 0.68 2.02 2.24 ;
        RECT  1.80 1.96 2.08 2.24 ;
        RECT  2.36 0.76 2.64 1.04 ;
        RECT  2.94 0.96 3.22 1.24 ;
        RECT  2.40 1.46 3.10 1.62 ;
        RECT  2.94 0.96 3.10 2.12 ;
        RECT  2.40 0.76 2.56 2.24 ;
        RECT  2.94 1.84 3.22 2.12 ;
        RECT  2.32 1.96 2.60 2.24 ;
        RECT  1.28 0.68 1.56 0.96 ;
        RECT  1.34 0.68 1.50 2.24 ;
        RECT  1.28 1.96 1.56 2.24 ;
        RECT  1.40 1.96 1.56 2.56 ;
        RECT  3.12 2.28 3.40 2.56 ;
        RECT  1.40 2.40 3.40 2.56 ;
    END
END XNR2SP4V1_0

MACRO XNR2SP2V1_0
    CLASS CORE ;
    FOREIGN XNR2SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 8.00  LAYER ME1  ;
        ANTENNADIFFAREA 3.69  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.31  LAYER ME1  ;
        ANTENNAMAXAREACAR 25.63  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.02 1.84 4.30 2.12 ;
        RECT  4.02 0.96 4.30 1.24 ;
        RECT  4.12 0.96 4.28 2.12 ;
        END
    END OUT
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.90 1.33 1.18 1.75 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.42 1.12 0.74 1.54 ;
        END
    END IN2
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.40 3.48 ;
        RECT  3.94 2.88 4.22 3.48 ;
        RECT  3.50 1.84 3.78 2.12 ;
        RECT  3.56 1.84 3.72 3.48 ;
        RECT  0.76 1.96 1.04 2.24 ;
        RECT  0.82 1.96 0.98 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.40 0.28 ;
        RECT  3.94 -0.28 4.22 0.32 ;
        RECT  3.50 0.64 3.78 0.92 ;
        RECT  3.56 -0.28 3.72 0.92 ;
        RECT  0.76 0.68 1.04 0.96 ;
        RECT  0.82 -0.28 0.98 0.96 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.68 0.52 0.96 ;
        RECT  0.10 1.96 0.52 2.24 ;
        RECT  0.10 0.68 0.26 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  1.92 0.44 3.08 0.60 ;
        RECT  2.80 0.44 3.08 0.72 ;
        RECT  1.92 0.44 2.08 0.96 ;
        RECT  1.80 0.68 2.08 0.96 ;
        RECT  1.86 0.68 2.02 2.24 ;
        RECT  1.80 1.96 2.08 2.24 ;
        RECT  2.36 0.76 2.64 1.04 ;
        RECT  2.94 0.96 3.22 1.24 ;
        RECT  2.40 1.46 3.10 1.62 ;
        RECT  2.94 0.96 3.10 2.12 ;
        RECT  2.40 0.76 2.56 2.24 ;
        RECT  2.94 1.84 3.22 2.12 ;
        RECT  2.32 1.96 2.60 2.24 ;
        RECT  1.28 0.68 1.56 0.96 ;
        RECT  1.34 0.68 1.50 2.24 ;
        RECT  1.28 1.96 1.56 2.24 ;
        RECT  1.40 1.96 1.56 2.56 ;
        RECT  3.12 2.28 3.40 2.56 ;
        RECT  1.40 2.40 3.40 2.56 ;
    END
END XNR2SP2V1_0

MACRO XNR2SP1V1_0
    CLASS CORE ;
    FOREIGN XNR2SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.42 1.12 0.74 1.54 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.90 1.33 1.18 1.75 ;
        END
    END IN1
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 8.05  LAYER ME1  ;
        ANTENNADIFFAREA 3.23  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.24  LAYER ME1  ;
        ANTENNAMAXAREACAR 34.22  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.98 1.84 4.28 2.12 ;
        RECT  4.12 0.96 4.28 2.12 ;
        RECT  3.98 0.96 4.28 1.24 ;
        END
    END OUT
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.40 0.28 ;
        RECT  3.94 -0.28 4.22 0.32 ;
        RECT  3.46 0.96 3.74 1.24 ;
        RECT  3.52 -0.28 3.68 1.24 ;
        RECT  0.76 0.68 1.04 0.96 ;
        RECT  0.82 -0.28 0.98 0.96 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.40 3.48 ;
        RECT  3.94 2.88 4.22 3.48 ;
        RECT  3.46 1.84 3.74 2.12 ;
        RECT  3.56 1.84 3.72 3.48 ;
        RECT  0.76 1.96 1.04 2.24 ;
        RECT  0.82 1.96 0.98 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.68 0.52 0.96 ;
        RECT  0.10 1.96 0.52 2.24 ;
        RECT  0.10 0.68 0.26 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  1.92 0.44 3.08 0.60 ;
        RECT  2.80 0.44 3.08 0.72 ;
        RECT  1.92 0.44 2.08 0.96 ;
        RECT  1.80 0.68 2.08 0.96 ;
        RECT  1.86 0.68 2.02 2.24 ;
        RECT  1.80 1.96 2.08 2.24 ;
        RECT  2.36 0.76 2.64 1.04 ;
        RECT  2.94 0.96 3.22 1.24 ;
        RECT  2.40 1.46 3.10 1.62 ;
        RECT  2.94 0.96 3.10 2.12 ;
        RECT  2.40 0.76 2.56 2.24 ;
        RECT  2.94 1.84 3.22 2.12 ;
        RECT  2.32 1.96 2.60 2.24 ;
        RECT  1.28 0.68 1.56 0.96 ;
        RECT  1.34 0.68 1.50 2.24 ;
        RECT  1.28 1.96 1.56 2.24 ;
        RECT  1.40 1.96 1.56 2.56 ;
        RECT  3.12 2.28 3.40 2.56 ;
        RECT  1.40 2.40 3.40 2.56 ;
    END
END XNR2SP1V1_0

MACRO TIE1SP8V1_0
    CLASS CORE ;
    FOREIGN TIE1SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 2.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 2.04  LAYER ME1  ;
        ANTENNADIFFAREA 1.64  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.66 1.84 1.94 2.12 ;
        RECT  0.62 1.84 1.94 2.00 ;
        RECT  0.62 1.84 0.90 2.12 ;
        RECT  0.62 1.46 0.78 2.12 ;
        RECT  0.46 1.46 0.78 1.74 ;
        END
    END OUT
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 2.80 0.28 ;
        RECT  2.24 -0.28 2.62 0.32 ;
        RECT  2.18 0.64 2.46 0.92 ;
        RECT  2.24 -0.28 2.40 0.92 ;
        RECT  1.14 0.64 1.42 0.92 ;
        RECT  1.20 -0.28 1.36 0.92 ;
        RECT  0.10 0.64 0.38 1.24 ;
        RECT  0.16 -0.28 0.32 1.24 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 2.80 3.48 ;
        RECT  2.24 2.88 2.62 3.48 ;
        RECT  2.18 2.16 2.46 2.44 ;
        RECT  2.24 2.16 2.40 3.48 ;
        RECT  1.14 2.16 1.42 2.44 ;
        RECT  1.20 2.16 1.36 3.48 ;
        RECT  0.10 2.16 0.38 2.44 ;
        RECT  0.16 2.16 0.32 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.64 0.90 1.24 ;
        RECT  1.66 0.96 1.94 1.24 ;
        RECT  0.62 1.08 1.94 1.24 ;
        RECT  1.78 0.96 1.94 1.56 ;
        RECT  1.78 1.40 2.28 1.56 ;
        RECT  2.00 1.40 2.28 1.68 ;
    END
END TIE1SP8V1_0

MACRO TIE1SP4V1_0
    CLASS CORE ;
    FOREIGN TIE1SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 1.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 1.21  LAYER ME1  ;
        ANTENNADIFFAREA 0.97  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.62 1.84 0.90 2.12 ;
        RECT  0.62 1.46 0.78 2.12 ;
        RECT  0.46 1.46 0.78 1.74 ;
        END
    END OUT
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 1.60 0.28 ;
        RECT  1.14 0.64 1.42 0.92 ;
        RECT  1.14 -0.28 1.42 0.32 ;
        RECT  1.20 -0.28 1.36 0.92 ;
        RECT  0.10 0.64 0.38 1.24 ;
        RECT  0.16 -0.28 0.32 1.24 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 1.60 3.48 ;
        RECT  1.14 2.88 1.42 3.48 ;
        RECT  1.14 2.16 1.42 2.44 ;
        RECT  1.20 2.16 1.36 3.48 ;
        RECT  0.10 2.16 0.38 2.44 ;
        RECT  0.16 2.16 0.32 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.64 0.90 1.24 ;
        RECT  0.62 1.08 1.12 1.24 ;
        RECT  0.96 1.08 1.12 1.68 ;
        RECT  0.96 1.40 1.24 1.68 ;
    END
END TIE1SP4V1_0

MACRO TIE1SP2V1_0
    CLASS CORE ;
    FOREIGN TIE1SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 1.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 0.83  LAYER ME1  ;
        ANTENNADIFFAREA 0.67  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.84 0.38 2.12 ;
        RECT  0.10 1.46 0.34 2.12 ;
        RECT  0.08 1.46 0.34 1.74 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 1.20 3.48 ;
        RECT  0.68 2.88 1.02 3.48 ;
        RECT  0.62 2.16 0.90 2.44 ;
        RECT  0.68 2.16 0.84 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 1.20 0.28 ;
        RECT  0.74 -0.28 1.02 0.32 ;
        RECT  0.10 0.64 0.38 1.24 ;
        RECT  0.16 -0.28 0.32 1.24 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.64 0.90 1.62 ;
    END
END TIE1SP2V1_0

MACRO TIE1SP1V1_0
    CLASS CORE ;
    FOREIGN TIE1SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 1.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 0.89  LAYER ME1  ;
        ANTENNADIFFAREA 0.45  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.84 0.38 2.12 ;
        RECT  0.10 1.46 0.34 2.12 ;
        RECT  0.08 1.46 0.34 1.74 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 1.20 3.48 ;
        RECT  0.68 2.88 1.02 3.48 ;
        RECT  0.62 1.84 0.90 2.12 ;
        RECT  0.68 1.84 0.84 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 1.20 0.28 ;
        RECT  0.74 -0.28 1.02 0.32 ;
        RECT  0.10 0.96 0.38 1.24 ;
        RECT  0.16 -0.28 0.32 1.24 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.96 0.90 1.62 ;
    END
END TIE1SP1V1_0

MACRO TIE0SP8V1_0
    CLASS CORE ;
    FOREIGN TIE0SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 2.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 2.25  LAYER ME1  ;
        ANTENNADIFFAREA 1.64  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.66 0.64 1.94 1.24 ;
        RECT  0.74 1.40 1.82 1.56 ;
        RECT  1.66 0.64 1.82 1.56 ;
        RECT  0.86 1.40 1.14 1.74 ;
        RECT  0.74 0.64 0.90 1.56 ;
        RECT  0.62 0.64 0.90 1.24 ;
        END
    END OUT
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 2.80 0.28 ;
        RECT  2.24 -0.28 2.62 0.32 ;
        RECT  2.18 0.64 2.46 1.24 ;
        RECT  2.24 -0.28 2.40 1.24 ;
        RECT  1.14 0.64 1.42 1.24 ;
        RECT  1.20 -0.28 1.36 1.24 ;
        RECT  0.10 0.64 0.38 1.24 ;
        RECT  0.16 -0.28 0.32 1.24 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 2.80 3.48 ;
        RECT  2.24 2.88 2.62 3.48 ;
        RECT  2.18 2.22 2.46 2.50 ;
        RECT  2.24 2.22 2.40 3.48 ;
        RECT  1.14 2.22 1.42 2.50 ;
        RECT  1.20 2.22 1.36 3.48 ;
        RECT  0.10 2.22 0.38 2.50 ;
        RECT  0.16 2.22 0.32 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  2.00 1.52 2.28 1.80 ;
        RECT  2.00 1.52 2.16 2.06 ;
        RECT  0.62 1.90 2.16 2.06 ;
        RECT  0.62 1.90 0.90 2.18 ;
        RECT  1.66 1.90 1.94 2.18 ;
    END
END TIE0SP8V1_0

MACRO TIE0SP4V1_0
    CLASS CORE ;
    FOREIGN TIE0SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 1.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 1.35  LAYER ME1  ;
        ANTENNADIFFAREA 0.97  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.62 0.64 0.90 1.24 ;
        RECT  0.46 1.46 0.78 1.74 ;
        RECT  0.62 0.64 0.78 1.74 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 1.60 3.48 ;
        RECT  1.14 2.88 1.42 3.48 ;
        RECT  1.14 2.22 1.42 2.50 ;
        RECT  1.20 2.22 1.36 3.48 ;
        RECT  0.10 2.22 0.38 2.50 ;
        RECT  0.16 2.22 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 1.60 0.28 ;
        RECT  1.14 0.64 1.42 1.24 ;
        RECT  1.14 -0.28 1.42 0.32 ;
        RECT  1.20 -0.28 1.36 1.24 ;
        RECT  0.10 0.64 0.38 1.24 ;
        RECT  0.16 -0.28 0.32 1.24 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.96 1.46 1.24 1.74 ;
        RECT  0.96 1.46 1.12 2.06 ;
        RECT  0.62 1.90 1.12 2.06 ;
        RECT  0.62 1.90 0.90 2.18 ;
    END
END TIE0SP4V1_0

MACRO TIE0SP2V1_0
    CLASS CORE ;
    FOREIGN TIE0SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 1.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 0.90  LAYER ME1  ;
        ANTENNADIFFAREA 0.67  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.20 0.64 0.48 1.24 ;
        RECT  0.08 1.46 0.36 1.74 ;
        RECT  0.20 0.64 0.36 1.74 ;
        END
    END OUT
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 1.20 0.28 ;
        RECT  0.74 -0.28 1.02 0.32 ;
        RECT  0.72 0.64 1.00 1.24 ;
        RECT  0.78 -0.28 0.94 1.24 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 1.20 3.48 ;
        RECT  0.74 2.88 1.02 3.48 ;
        RECT  0.20 2.16 0.48 2.44 ;
        RECT  0.26 2.16 0.42 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.74 1.40 1.02 1.68 ;
        RECT  0.78 1.40 0.94 2.12 ;
        RECT  0.72 1.84 1.00 2.12 ;
    END
END TIE0SP2V1_0

MACRO TIE0SP1V1_0
    CLASS CORE ;
    FOREIGN TIE0SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 1.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 0.86  LAYER ME1  ;
        ANTENNADIFFAREA 0.45  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.20 0.96 0.48 1.24 ;
        RECT  0.08 1.46 0.36 1.74 ;
        RECT  0.20 0.96 0.36 1.74 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 1.20 3.48 ;
        RECT  0.74 2.88 1.02 3.48 ;
        RECT  0.20 1.90 0.48 2.18 ;
        RECT  0.26 1.90 0.42 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 1.20 0.28 ;
        RECT  0.74 -0.28 1.02 0.32 ;
        RECT  0.72 0.96 1.00 1.24 ;
        RECT  0.78 -0.28 0.94 1.24 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.74 1.40 1.02 1.68 ;
        RECT  0.78 1.40 0.94 2.18 ;
        RECT  0.72 1.90 1.00 2.18 ;
    END
END TIE0SP1V1_0

MACRO OR3SP8V1_0
    CLASS CORE ;
    FOREIGN OR3SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.46 1.62 1.86 ;
        END
    END IN3
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 7.97  LAYER ME1  ;
        ANTENNADIFFAREA 4.62  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.58  LAYER ME1  ;
        ANTENNAMAXAREACAR 13.84  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.24 0.70 3.54 0.98 ;
        RECT  3.12 2.06 3.40 2.66 ;
        RECT  3.24 0.70 3.40 2.66 ;
        RECT  2.26 1.52 3.40 1.68 ;
        RECT  2.22 0.70 2.50 0.98 ;
        RECT  2.08 2.06 2.42 2.66 ;
        RECT  2.26 0.70 2.42 2.66 ;
        END
    END OUT
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.46 0.38 1.86 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.46 1.14 1.86 ;
        END
    END IN2
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.40 3.48 ;
        RECT  3.70 2.88 4.22 3.48 ;
        RECT  3.64 2.06 3.92 2.66 ;
        RECT  3.70 2.06 3.86 3.48 ;
        RECT  2.60 2.06 2.88 2.66 ;
        RECT  2.66 2.06 2.82 3.48 ;
        RECT  1.56 2.06 1.84 2.66 ;
        RECT  1.62 2.06 1.78 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.40 0.28 ;
        RECT  3.84 -0.28 4.22 0.32 ;
        RECT  3.78 0.58 4.06 0.86 ;
        RECT  3.84 -0.28 4.00 0.86 ;
        RECT  2.74 0.58 3.02 0.86 ;
        RECT  2.80 -0.28 2.96 0.86 ;
        RECT  1.70 0.58 1.98 0.86 ;
        RECT  1.76 -0.28 1.92 0.86 ;
        RECT  0.62 0.64 0.90 0.92 ;
        RECT  0.68 -0.28 0.84 0.92 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.64 0.38 0.92 ;
        RECT  1.14 0.64 1.42 0.92 ;
        RECT  0.22 0.64 0.38 1.30 ;
        RECT  1.14 0.64 1.30 1.30 ;
        RECT  0.22 1.14 2.10 1.30 ;
        RECT  1.82 1.14 2.10 1.56 ;
        RECT  0.54 1.14 0.70 2.44 ;
        RECT  0.24 2.16 0.70 2.44 ;
    END
END OR3SP8V1_0

MACRO OR3SP4V1_0
    CLASS CORE ;
    FOREIGN OR3SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.46 1.14 1.86 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.46 1.62 1.86 ;
        END
    END IN3
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.46 0.38 1.86 ;
        END
    END IN1
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 5.27  LAYER ME1  ;
        ANTENNADIFFAREA 3.07  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.29  LAYER ME1  ;
        ANTENNAMAXAREACAR 18.31  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.26 1.52 2.68 1.68 ;
        RECT  2.22 0.70 2.50 0.98 ;
        RECT  2.08 2.06 2.42 2.66 ;
        RECT  2.26 0.70 2.42 2.66 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 3.20 3.48 ;
        RECT  2.66 2.88 3.02 3.48 ;
        RECT  2.60 2.06 2.88 2.66 ;
        RECT  2.66 2.06 2.82 3.48 ;
        RECT  1.56 2.06 1.84 2.66 ;
        RECT  1.62 2.06 1.78 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 3.20 0.28 ;
        RECT  2.74 0.58 3.02 0.86 ;
        RECT  2.74 -0.28 3.02 0.32 ;
        RECT  2.80 -0.28 2.96 0.86 ;
        RECT  1.70 0.58 1.98 0.86 ;
        RECT  1.76 -0.28 1.92 0.86 ;
        RECT  0.62 0.64 0.90 0.92 ;
        RECT  0.68 -0.28 0.84 0.92 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.64 0.38 0.92 ;
        RECT  1.14 0.64 1.42 0.92 ;
        RECT  0.22 0.64 0.38 1.30 ;
        RECT  1.14 0.64 1.30 1.30 ;
        RECT  0.22 1.14 2.10 1.30 ;
        RECT  1.82 1.14 2.10 1.56 ;
        RECT  0.54 1.14 0.70 2.44 ;
        RECT  0.24 2.16 0.70 2.44 ;
    END
END OR3SP4V1_0

MACRO OR3SP2V1_0
    CLASS CORE ;
    FOREIGN OR3SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 2.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 4.53  LAYER ME1  ;
        ANTENNADIFFAREA 2.46  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.14  LAYER ME1  ;
        ANTENNAMAXAREACAR 31.44  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.08 2.06 2.68 2.22 ;
        RECT  2.52 0.80 2.68 2.22 ;
        RECT  2.22 0.80 2.68 0.96 ;
        RECT  2.22 0.68 2.50 0.96 ;
        RECT  2.08 2.06 2.36 2.66 ;
        END
    END OUT
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.44 0.38 1.86 ;
        END
    END IN1
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.34 1.46 1.92 1.74 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.44 1.14 1.86 ;
        END
    END IN2
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 2.80 0.28 ;
        RECT  2.34 -0.28 2.62 0.32 ;
        RECT  1.70 0.54 1.98 0.82 ;
        RECT  1.76 -0.28 1.92 0.82 ;
        RECT  0.62 0.64 0.90 0.92 ;
        RECT  0.68 -0.28 0.84 0.92 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 2.80 3.48 ;
        RECT  2.34 2.88 2.62 3.48 ;
        RECT  1.56 2.06 1.84 2.66 ;
        RECT  1.62 2.06 1.78 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.64 0.38 0.92 ;
        RECT  1.14 0.64 1.42 0.92 ;
        RECT  0.22 0.64 0.38 1.28 ;
        RECT  1.14 0.64 1.30 1.28 ;
        RECT  0.22 1.12 2.24 1.28 ;
        RECT  2.08 1.12 2.24 1.63 ;
        RECT  2.08 1.35 2.36 1.63 ;
        RECT  0.54 1.12 0.70 2.44 ;
        RECT  0.24 2.16 0.70 2.44 ;
    END
END OR3SP2V1_0

MACRO OR3SP1V1_0
    CLASS CORE ;
    FOREIGN OR3SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 2.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 4.45  LAYER ME1  ;
        ANTENNADIFFAREA 2.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 66.23  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.04 2.16 2.68 2.32 ;
        RECT  2.52 0.76 2.68 2.32 ;
        RECT  2.18 0.76 2.68 0.92 ;
        RECT  2.18 0.64 2.46 0.92 ;
        RECT  2.04 2.16 2.32 2.44 ;
        END
    END OUT
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.34 1.46 1.94 1.74 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.44 1.14 1.86 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.44 0.38 1.86 ;
        END
    END IN1
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 2.80 0.28 ;
        RECT  2.34 -0.28 2.62 0.32 ;
        RECT  1.66 0.64 1.94 0.92 ;
        RECT  1.72 -0.28 1.88 0.92 ;
        RECT  0.62 0.64 0.90 0.92 ;
        RECT  0.68 -0.28 0.84 0.92 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 2.80 3.48 ;
        RECT  2.34 2.88 2.62 3.48 ;
        RECT  1.52 2.16 1.80 2.44 ;
        RECT  1.58 2.16 1.74 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.64 0.38 0.92 ;
        RECT  1.14 0.64 1.42 0.92 ;
        RECT  0.22 0.64 0.38 1.28 ;
        RECT  1.14 0.64 1.30 1.28 ;
        RECT  0.22 1.12 2.35 1.28 ;
        RECT  2.07 1.08 2.35 1.36 ;
        RECT  0.54 1.12 0.70 2.44 ;
        RECT  0.24 2.16 0.70 2.44 ;
    END
END OR3SP1V1_0

MACRO OR3NAND2SP8V1_0
    CLASS CORE ;
    FOREIGN OR3NAND2SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 11.96  LAYER ME1  ;
        ANTENNADIFFAREA 6.59  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.71  LAYER ME1  ;
        ANTENNAMAXAREACAR 16.84  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.30 1.98 5.58 2.58 ;
        RECT  5.30 0.64 5.58 1.24 ;
        RECT  5.30 0.64 5.46 2.58 ;
        RECT  4.34 1.52 5.46 1.68 ;
        RECT  4.34 1.46 4.74 1.74 ;
        RECT  4.26 1.98 4.54 2.58 ;
        RECT  4.26 0.64 4.54 1.24 ;
        RECT  4.34 0.64 4.50 2.58 ;
        END
    END OUT
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.00 1.40 2.28 1.82 ;
        END
    END IN4
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.40 0.70 1.82 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.40 1.16 1.82 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.32 1.40 1.64 1.82 ;
        END
    END IN3
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 6.40 0.28 ;
        RECT  5.88 -0.28 6.22 0.32 ;
        RECT  5.82 0.64 6.10 1.24 ;
        RECT  5.88 -0.28 6.04 1.24 ;
        RECT  4.78 0.64 5.06 1.24 ;
        RECT  4.84 -0.28 5.00 1.24 ;
        RECT  3.74 0.64 4.02 1.24 ;
        RECT  3.80 -0.28 3.96 1.24 ;
        RECT  2.66 0.64 2.94 0.92 ;
        RECT  2.72 -0.28 2.88 0.92 ;
        RECT  1.66 0.64 1.94 0.92 ;
        RECT  1.72 -0.28 1.88 0.92 ;
        RECT  0.62 0.64 0.90 0.92 ;
        RECT  0.68 -0.28 0.84 0.92 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 6.40 3.48 ;
        RECT  5.88 2.88 6.22 3.48 ;
        RECT  5.82 1.98 6.10 2.58 ;
        RECT  5.88 1.98 6.04 3.48 ;
        RECT  4.78 1.98 5.06 2.58 ;
        RECT  4.84 1.98 5.00 3.48 ;
        RECT  3.74 1.98 4.02 2.58 ;
        RECT  3.80 1.98 3.96 3.48 ;
        RECT  1.52 2.02 1.80 2.30 ;
        RECT  1.58 2.02 1.74 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.08 0.64 0.38 0.92 ;
        RECT  1.14 0.64 1.42 0.92 ;
        RECT  1.14 0.64 1.30 1.24 ;
        RECT  0.08 1.08 1.30 1.24 ;
        RECT  0.08 2.02 0.52 2.30 ;
        RECT  0.08 0.64 0.24 2.76 ;
        RECT  0.08 2.48 0.38 2.76 ;
        RECT  2.18 0.64 2.46 0.92 ;
        RECT  2.30 0.64 2.46 1.24 ;
        RECT  2.44 1.46 2.76 1.74 ;
        RECT  2.44 1.08 2.60 2.30 ;
        RECT  2.04 2.02 2.60 2.30 ;
        RECT  3.18 0.64 3.46 0.92 ;
        RECT  3.24 1.52 4.16 1.68 ;
        RECT  3.88 1.46 4.16 1.74 ;
        RECT  3.24 0.64 3.40 2.18 ;
        RECT  2.80 2.02 3.40 2.18 ;
        RECT  2.80 2.02 3.08 2.30 ;
    END
END OR3NAND2SP8V1_0

MACRO OR3NAND2SP4V1_0
    CLASS CORE ;
    FOREIGN OR3NAND2SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.32 1.40 1.64 1.82 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.40 1.16 1.82 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.40 0.70 1.82 ;
        END
    END IN1
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.00 1.40 2.28 1.82 ;
        END
    END IN4
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 9.62  LAYER ME1  ;
        ANTENNADIFFAREA 4.77  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.42  LAYER ME1  ;
        ANTENNAMAXAREACAR 22.78  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.34 1.46 4.74 1.74 ;
        RECT  4.26 1.98 4.54 2.58 ;
        RECT  4.26 0.64 4.54 1.24 ;
        RECT  4.34 0.64 4.50 2.58 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 5.20 3.48 ;
        RECT  4.78 1.98 5.06 2.58 ;
        RECT  4.74 2.88 5.02 3.48 ;
        RECT  4.84 1.98 5.00 3.48 ;
        RECT  3.74 1.98 4.02 2.58 ;
        RECT  3.80 1.98 3.96 3.48 ;
        RECT  1.52 2.02 1.80 2.30 ;
        RECT  1.58 2.02 1.74 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 5.20 0.28 ;
        RECT  4.78 0.64 5.06 1.24 ;
        RECT  4.74 -0.28 5.02 0.32 ;
        RECT  4.84 -0.28 5.00 1.24 ;
        RECT  3.74 0.64 4.02 1.24 ;
        RECT  3.80 -0.28 3.96 1.24 ;
        RECT  2.66 0.64 2.94 0.92 ;
        RECT  2.72 -0.28 2.88 0.92 ;
        RECT  1.66 0.64 1.94 0.92 ;
        RECT  1.72 -0.28 1.88 0.92 ;
        RECT  0.62 0.64 0.90 0.92 ;
        RECT  0.68 -0.28 0.84 0.92 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.08 0.64 0.38 0.92 ;
        RECT  1.14 0.64 1.42 0.92 ;
        RECT  1.14 0.64 1.30 1.24 ;
        RECT  0.08 1.08 1.30 1.24 ;
        RECT  0.08 2.02 0.52 2.30 ;
        RECT  0.08 0.64 0.24 2.76 ;
        RECT  0.08 2.48 0.38 2.76 ;
        RECT  2.18 0.64 2.46 0.92 ;
        RECT  2.30 0.64 2.46 1.24 ;
        RECT  2.44 1.46 2.76 1.74 ;
        RECT  2.44 1.08 2.60 2.30 ;
        RECT  2.04 2.02 2.60 2.30 ;
        RECT  3.18 0.64 3.46 0.92 ;
        RECT  3.24 1.52 4.16 1.68 ;
        RECT  3.88 1.46 4.16 1.74 ;
        RECT  3.24 0.64 3.40 2.18 ;
        RECT  2.80 2.02 3.40 2.18 ;
        RECT  2.80 2.02 3.08 2.30 ;
    END
END OR3NAND2SP4V1_0

MACRO OR3NAND2SP2V1_0
    CLASS CORE ;
    FOREIGN OR3NAND2SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 8.74  LAYER ME1  ;
        ANTENNADIFFAREA 4.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.28  LAYER ME1  ;
        ANTENNAMAXAREACAR 31.38  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.34 1.46 4.72 1.74 ;
        RECT  4.26 1.98 4.54 2.58 ;
        RECT  4.26 0.64 4.54 1.24 ;
        RECT  4.34 0.64 4.50 2.58 ;
        END
    END OUT
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.00 1.40 2.28 1.82 ;
        END
    END IN4
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.40 0.70 1.82 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.40 1.16 1.82 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.32 1.40 1.64 1.82 ;
        END
    END IN3
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.80 0.28 ;
        RECT  4.34 -0.28 4.62 0.32 ;
        RECT  3.74 0.64 4.02 1.24 ;
        RECT  3.80 -0.28 3.96 1.24 ;
        RECT  2.66 0.64 2.94 0.92 ;
        RECT  2.72 -0.28 2.88 0.92 ;
        RECT  1.66 0.64 1.94 0.92 ;
        RECT  1.72 -0.28 1.88 0.92 ;
        RECT  0.62 0.64 0.90 0.92 ;
        RECT  0.68 -0.28 0.84 0.92 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.80 3.48 ;
        RECT  4.34 2.88 4.62 3.48 ;
        RECT  3.74 1.98 4.02 2.58 ;
        RECT  3.80 1.98 3.96 3.48 ;
        RECT  1.52 2.02 1.80 2.30 ;
        RECT  1.58 2.02 1.74 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.08 0.64 0.38 0.92 ;
        RECT  1.14 0.64 1.42 0.92 ;
        RECT  1.14 0.64 1.30 1.24 ;
        RECT  0.08 1.08 1.30 1.24 ;
        RECT  0.08 2.02 0.52 2.30 ;
        RECT  0.08 0.64 0.24 2.76 ;
        RECT  0.08 2.48 0.38 2.76 ;
        RECT  2.18 0.64 2.46 0.92 ;
        RECT  2.30 0.64 2.46 1.24 ;
        RECT  2.44 1.46 2.76 1.74 ;
        RECT  2.44 1.08 2.60 2.30 ;
        RECT  2.04 2.02 2.60 2.30 ;
        RECT  3.18 0.64 3.46 0.92 ;
        RECT  3.24 1.52 4.16 1.68 ;
        RECT  3.88 1.46 4.16 1.74 ;
        RECT  3.24 0.64 3.40 2.18 ;
        RECT  2.80 2.02 3.40 2.18 ;
        RECT  2.80 2.02 3.08 2.30 ;
    END
END OR3NAND2SP2V1_0

MACRO OR3NAND2SP1V1_0
    CLASS CORE ;
    FOREIGN OR3NAND2SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 8.08  LAYER ME1  ;
        ANTENNADIFFAREA 3.55  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        ANTENNAMAXAREACAR 40.10  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.34 1.46 4.72 1.74 ;
        RECT  4.22 2.02 4.50 2.30 ;
        RECT  4.34 0.64 4.50 2.30 ;
        RECT  4.22 0.64 4.50 0.92 ;
        END
    END OUT
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.32 1.40 1.64 1.82 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.40 1.16 1.82 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.40 0.70 1.82 ;
        END
    END IN1
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.00 1.40 2.28 1.82 ;
        END
    END IN4
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.80 0.28 ;
        RECT  4.34 -0.28 4.62 0.32 ;
        RECT  3.70 0.64 3.98 0.92 ;
        RECT  3.76 -0.28 3.92 0.92 ;
        RECT  2.66 0.64 2.94 0.92 ;
        RECT  2.72 -0.28 2.88 0.92 ;
        RECT  1.66 0.64 1.94 0.92 ;
        RECT  1.72 -0.28 1.88 0.92 ;
        RECT  0.62 0.64 0.90 0.92 ;
        RECT  0.68 -0.28 0.84 0.92 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.80 3.48 ;
        RECT  4.34 2.88 4.62 3.48 ;
        RECT  3.70 2.02 3.98 2.30 ;
        RECT  3.76 2.02 3.92 3.48 ;
        RECT  1.52 2.02 1.80 2.30 ;
        RECT  1.58 2.02 1.74 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.08 0.64 0.38 0.92 ;
        RECT  1.14 0.64 1.42 0.92 ;
        RECT  1.14 0.64 1.30 1.24 ;
        RECT  0.08 1.08 1.30 1.24 ;
        RECT  0.08 2.02 0.52 2.30 ;
        RECT  0.08 0.64 0.24 2.76 ;
        RECT  0.08 2.48 0.38 2.76 ;
        RECT  2.18 0.64 2.46 0.92 ;
        RECT  2.30 0.64 2.46 1.24 ;
        RECT  2.44 1.46 2.76 1.74 ;
        RECT  2.44 1.08 2.60 2.30 ;
        RECT  2.04 2.02 2.60 2.30 ;
        RECT  3.18 0.64 3.46 0.92 ;
        RECT  3.24 1.52 4.16 1.68 ;
        RECT  3.88 1.46 4.16 1.74 ;
        RECT  3.24 0.64 3.40 2.18 ;
        RECT  2.80 2.02 3.40 2.18 ;
        RECT  2.80 2.02 3.08 2.30 ;
    END
END OR3NAND2SP1V1_0

MACRO OR3I2SP8V1_0
    CLASS CORE ;
    FOREIGN OR3I2SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 11.07  LAYER ME1  ;
        ANTENNADIFFAREA 5.53  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.71  LAYER ME1  ;
        ANTENNAMAXAREACAR 15.58  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.88 1.04 5.20 1.20 ;
        RECT  4.92 0.60 5.20 1.20 ;
        RECT  4.78 2.06 5.06 2.66 ;
        RECT  3.74 2.06 5.06 2.22 ;
        RECT  4.12 1.04 4.28 2.22 ;
        RECT  3.88 0.60 4.16 1.20 ;
        RECT  3.74 2.06 4.02 2.66 ;
        END
    END OUT
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.86 1.46 3.26 1.74 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.42 1.39 0.70 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.18 1.81 ;
        END
    END IN1
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 6.00 0.28 ;
        RECT  5.50 -0.28 5.82 0.32 ;
        RECT  5.44 0.60 5.72 1.20 ;
        RECT  5.50 -0.28 5.66 1.20 ;
        RECT  4.40 0.60 4.68 0.88 ;
        RECT  4.46 -0.28 4.62 0.88 ;
        RECT  3.36 0.60 3.64 0.88 ;
        RECT  3.42 -0.28 3.58 0.88 ;
        RECT  2.28 0.64 2.56 0.92 ;
        RECT  2.34 -0.28 2.50 0.92 ;
        RECT  0.76 0.64 1.04 0.92 ;
        RECT  0.82 -0.28 0.98 0.92 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 6.00 3.48 ;
        RECT  5.38 2.88 5.82 3.48 ;
        RECT  5.30 2.06 5.58 2.66 ;
        RECT  5.38 2.06 5.54 3.48 ;
        RECT  4.26 2.38 4.54 2.66 ;
        RECT  4.32 2.38 4.48 3.48 ;
        RECT  3.22 2.06 3.50 2.66 ;
        RECT  3.28 2.06 3.44 3.48 ;
        RECT  0.76 1.97 1.04 2.25 ;
        RECT  0.82 1.97 0.98 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.64 0.52 0.92 ;
        RECT  0.10 1.97 0.52 2.25 ;
        RECT  0.10 0.64 0.26 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  1.28 0.64 1.60 0.92 ;
        RECT  1.44 1.46 1.88 1.74 ;
        RECT  1.44 0.64 1.60 2.25 ;
        RECT  1.28 1.97 1.60 2.25 ;
        RECT  1.76 0.64 2.04 0.92 ;
        RECT  2.80 0.64 3.08 0.92 ;
        RECT  1.88 0.64 2.04 1.28 ;
        RECT  2.80 0.64 2.96 1.28 ;
        RECT  1.88 1.12 3.62 1.28 ;
        RECT  3.46 1.12 3.62 1.64 ;
        RECT  3.46 1.36 3.74 1.64 ;
        RECT  2.06 1.12 2.22 2.44 ;
        RECT  1.90 2.16 2.36 2.44 ;
    END
END OR3I2SP8V1_0

MACRO OR3I2SP4V1_0
    CLASS CORE ;
    FOREIGN OR3I2SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.18 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.42 1.39 0.70 1.81 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.86 1.46 3.26 1.74 ;
        END
    END IN3
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 8.95  LAYER ME1  ;
        ANTENNADIFFAREA 4.19  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.42  LAYER ME1  ;
        ANTENNAMAXAREACAR 21.19  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.90 1.52 4.28 1.68 ;
        RECT  3.88 0.60 4.16 1.20 ;
        RECT  3.74 2.06 4.06 2.66 ;
        RECT  3.90 0.60 4.06 2.66 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.80 3.48 ;
        RECT  4.32 2.88 4.62 3.48 ;
        RECT  4.26 2.06 4.54 2.66 ;
        RECT  4.32 2.06 4.48 3.48 ;
        RECT  3.22 2.06 3.50 2.66 ;
        RECT  3.28 2.06 3.44 3.48 ;
        RECT  0.76 1.97 1.04 2.25 ;
        RECT  0.82 1.97 0.98 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.80 0.28 ;
        RECT  4.40 0.60 4.68 1.20 ;
        RECT  4.46 -0.28 4.62 1.20 ;
        RECT  4.34 -0.28 4.62 0.32 ;
        RECT  3.36 0.60 3.64 0.88 ;
        RECT  3.42 -0.28 3.58 0.88 ;
        RECT  2.28 0.64 2.56 0.92 ;
        RECT  2.34 -0.28 2.50 0.92 ;
        RECT  0.76 0.64 1.04 0.92 ;
        RECT  0.82 -0.28 0.98 0.92 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.64 0.52 0.92 ;
        RECT  0.10 1.97 0.52 2.25 ;
        RECT  0.10 0.64 0.26 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  1.28 0.64 1.60 0.92 ;
        RECT  1.44 1.46 1.88 1.74 ;
        RECT  1.44 0.64 1.60 2.25 ;
        RECT  1.28 1.97 1.60 2.25 ;
        RECT  1.76 0.64 2.04 0.92 ;
        RECT  2.80 0.64 3.08 0.92 ;
        RECT  1.88 0.64 2.04 1.28 ;
        RECT  2.80 0.64 2.96 1.28 ;
        RECT  1.88 1.12 3.62 1.28 ;
        RECT  3.46 1.12 3.62 1.64 ;
        RECT  3.46 1.36 3.74 1.64 ;
        RECT  2.06 1.12 2.22 2.44 ;
        RECT  1.90 2.16 2.36 2.44 ;
    END
END OR3I2SP4V1_0

MACRO OR3I2SP2V1_0
    CLASS CORE ;
    FOREIGN OR3I2SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 8.14  LAYER ME1  ;
        ANTENNADIFFAREA 3.58  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.28  LAYER ME1  ;
        ANTENNAMAXAREACAR 29.24  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.74 2.06 4.28 2.22 ;
        RECT  4.12 0.54 4.28 2.22 ;
        RECT  3.88 0.54 4.28 1.14 ;
        RECT  3.74 2.06 4.02 2.66 ;
        END
    END OUT
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.86 1.46 3.26 1.74 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.42 1.39 0.70 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.18 1.81 ;
        END
    END IN1
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.40 0.28 ;
        RECT  3.94 -0.28 4.22 0.32 ;
        RECT  3.36 0.54 3.64 0.82 ;
        RECT  3.42 -0.28 3.58 0.82 ;
        RECT  2.28 0.64 2.56 0.92 ;
        RECT  2.34 -0.28 2.50 0.92 ;
        RECT  0.76 0.64 1.04 0.92 ;
        RECT  0.82 -0.28 0.98 0.92 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.40 3.48 ;
        RECT  3.94 2.88 4.22 3.48 ;
        RECT  3.22 2.06 3.50 2.66 ;
        RECT  3.28 2.06 3.44 3.48 ;
        RECT  0.76 1.97 1.04 2.25 ;
        RECT  0.82 1.97 0.98 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.64 0.52 0.92 ;
        RECT  0.10 1.97 0.52 2.25 ;
        RECT  0.10 0.64 0.26 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  1.28 0.64 1.60 0.92 ;
        RECT  1.44 1.46 1.88 1.74 ;
        RECT  1.44 0.64 1.60 2.25 ;
        RECT  1.28 1.97 1.60 2.25 ;
        RECT  1.76 0.64 2.04 0.92 ;
        RECT  2.80 0.64 3.08 0.92 ;
        RECT  1.88 0.64 2.04 1.28 ;
        RECT  2.80 0.64 2.96 1.28 ;
        RECT  1.88 1.12 3.70 1.28 ;
        RECT  3.54 1.12 3.70 1.57 ;
        RECT  3.54 1.29 3.82 1.57 ;
        RECT  2.06 1.12 2.22 2.44 ;
        RECT  1.90 2.16 2.36 2.44 ;
    END
END OR3I2SP2V1_0

MACRO OR3I2SP1V1_0
    CLASS CORE ;
    FOREIGN OR3I2SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 7.90  LAYER ME1  ;
        ANTENNADIFFAREA 3.12  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        ANTENNAMAXAREACAR 39.21  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.70 2.16 4.28 2.32 ;
        RECT  4.12 0.76 4.28 2.32 ;
        RECT  3.84 0.64 4.12 0.92 ;
        RECT  3.70 2.16 3.98 2.44 ;
        END
    END OUT
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.86 1.46 3.26 1.74 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.42 1.39 0.70 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.18 1.81 ;
        END
    END IN1
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.40 0.28 ;
        RECT  3.94 -0.28 4.22 0.32 ;
        RECT  3.32 0.64 3.60 0.92 ;
        RECT  3.38 -0.28 3.54 0.92 ;
        RECT  2.28 0.64 2.56 0.92 ;
        RECT  2.34 -0.28 2.50 0.92 ;
        RECT  0.76 0.64 1.04 0.92 ;
        RECT  0.82 -0.28 0.98 0.92 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.40 3.48 ;
        RECT  3.94 2.88 4.22 3.48 ;
        RECT  3.18 2.16 3.46 2.44 ;
        RECT  3.24 2.16 3.40 3.48 ;
        RECT  0.76 1.97 1.04 2.25 ;
        RECT  0.82 1.97 0.98 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.64 0.52 0.92 ;
        RECT  0.10 1.97 0.52 2.25 ;
        RECT  0.10 0.64 0.26 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  1.28 0.64 1.60 0.92 ;
        RECT  1.44 1.46 1.88 1.74 ;
        RECT  1.44 0.64 1.60 2.25 ;
        RECT  1.28 1.97 1.60 2.25 ;
        RECT  1.76 0.64 2.04 0.92 ;
        RECT  2.80 0.64 3.08 0.92 ;
        RECT  1.88 0.64 2.04 1.28 ;
        RECT  2.80 0.64 2.96 1.28 ;
        RECT  1.88 1.12 3.81 1.28 ;
        RECT  3.53 1.08 3.81 1.36 ;
        RECT  2.06 1.12 2.22 2.44 ;
        RECT  1.90 2.16 2.36 2.44 ;
    END
END OR3I2SP1V1_0

MACRO OR3I1SP8V1_0
    CLASS CORE ;
    FOREIGN OR3I1SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 9.93  LAYER ME1  ;
        ANTENNADIFFAREA 5.26  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.64  LAYER ME1  ;
        ANTENNAMAXAREACAR 15.44  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.26 0.60 4.54 1.20 ;
        RECT  4.12 2.06 4.42 2.66 ;
        RECT  4.26 0.60 4.42 2.66 ;
        RECT  3.32 1.52 4.42 1.68 ;
        RECT  3.22 0.60 3.50 1.20 ;
        RECT  3.32 0.60 3.48 1.93 ;
        RECT  3.08 2.06 3.44 2.66 ;
        RECT  3.28 1.77 3.44 2.66 ;
        END
    END OUT
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.34 1.46 2.72 1.74 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.72 1.44 2.04 1.86 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 5.20 3.48 ;
        RECT  4.70 2.88 5.02 3.48 ;
        RECT  4.64 2.06 4.92 2.66 ;
        RECT  4.70 2.06 4.86 3.48 ;
        RECT  3.60 2.06 3.88 2.66 ;
        RECT  3.66 2.06 3.82 3.48 ;
        RECT  2.56 2.06 2.84 2.66 ;
        RECT  2.62 2.06 2.78 3.48 ;
        RECT  0.10 2.16 0.38 2.44 ;
        RECT  0.16 2.16 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 5.20 0.28 ;
        RECT  4.78 0.60 5.06 1.20 ;
        RECT  4.74 -0.28 5.02 0.32 ;
        RECT  4.84 -0.28 5.00 1.20 ;
        RECT  3.74 0.60 4.02 1.20 ;
        RECT  3.80 -0.28 3.96 1.20 ;
        RECT  2.70 0.60 2.98 0.88 ;
        RECT  2.76 -0.28 2.92 0.88 ;
        RECT  1.62 0.64 1.90 0.92 ;
        RECT  1.68 -0.28 1.84 0.92 ;
        RECT  0.10 0.64 0.38 0.92 ;
        RECT  0.16 -0.28 0.32 0.92 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.64 0.94 0.92 ;
        RECT  0.78 1.46 1.22 1.74 ;
        RECT  0.78 0.64 0.94 2.44 ;
        RECT  0.62 2.16 0.94 2.44 ;
        RECT  1.10 0.64 1.38 0.92 ;
        RECT  2.14 0.64 2.42 0.92 ;
        RECT  1.22 0.64 1.38 1.28 ;
        RECT  2.14 0.64 2.30 1.28 ;
        RECT  1.22 1.12 3.04 1.28 ;
        RECT  2.88 1.12 3.04 1.66 ;
        RECT  2.88 1.38 3.16 1.66 ;
        RECT  1.40 1.12 1.56 2.44 ;
        RECT  1.24 2.16 1.70 2.44 ;
    END
END OR3I1SP8V1_0

MACRO OR3I1SP4V1_0
    CLASS CORE ;
    FOREIGN OR3I1SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.72 1.44 2.04 1.86 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.34 1.46 2.72 1.74 ;
        END
    END IN3
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 8.01  LAYER ME1  ;
        ANTENNADIFFAREA 3.84  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.36  LAYER ME1  ;
        ANTENNAMAXAREACAR 22.55  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.22 0.60 3.50 1.20 ;
        RECT  3.32 0.60 3.48 1.93 ;
        RECT  3.08 2.06 3.44 2.66 ;
        RECT  3.28 1.77 3.44 2.66 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.40 3.48 ;
        RECT  3.66 2.88 4.22 3.48 ;
        RECT  3.60 2.06 3.88 2.66 ;
        RECT  3.66 2.06 3.82 3.48 ;
        RECT  2.56 2.06 2.84 2.66 ;
        RECT  2.62 2.06 2.78 3.48 ;
        RECT  0.10 2.16 0.38 2.44 ;
        RECT  0.16 2.16 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.40 0.28 ;
        RECT  3.80 -0.28 4.22 0.32 ;
        RECT  3.74 0.60 4.02 1.20 ;
        RECT  3.80 -0.28 3.96 1.20 ;
        RECT  2.70 0.60 2.98 0.88 ;
        RECT  2.76 -0.28 2.92 0.88 ;
        RECT  1.62 0.64 1.90 0.92 ;
        RECT  1.68 -0.28 1.84 0.92 ;
        RECT  0.10 0.64 0.38 0.92 ;
        RECT  0.16 -0.28 0.32 0.92 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.64 0.94 0.92 ;
        RECT  0.78 1.46 1.22 1.74 ;
        RECT  0.78 0.64 0.94 2.44 ;
        RECT  0.62 2.16 0.94 2.44 ;
        RECT  1.10 0.64 1.38 0.92 ;
        RECT  2.14 0.64 2.42 0.92 ;
        RECT  1.22 0.64 1.38 1.28 ;
        RECT  2.14 0.64 2.30 1.28 ;
        RECT  1.22 1.12 3.04 1.28 ;
        RECT  2.88 1.12 3.04 1.66 ;
        RECT  2.88 1.38 3.16 1.66 ;
        RECT  1.40 1.12 1.56 2.44 ;
        RECT  1.24 2.16 1.70 2.44 ;
    END
END OR3I1SP4V1_0

MACRO OR3I1SP2V1_0
    CLASS CORE ;
    FOREIGN OR3I1SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 6.71  LAYER ME1  ;
        ANTENNADIFFAREA 3.10  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.21  LAYER ME1  ;
        ANTENNAMAXAREACAR 31.78  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.22 0.60 3.50 1.20 ;
        RECT  3.08 2.06 3.48 2.66 ;
        RECT  3.32 0.60 3.48 2.66 ;
        END
    END OUT
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.34 1.46 2.72 1.74 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.72 1.44 2.04 1.86 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 3.60 0.28 ;
        RECT  3.14 -0.28 3.42 0.32 ;
        RECT  2.70 0.60 2.98 0.88 ;
        RECT  2.76 -0.28 2.92 0.88 ;
        RECT  1.62 0.64 1.90 0.92 ;
        RECT  1.68 -0.28 1.84 0.92 ;
        RECT  0.10 0.64 0.38 0.92 ;
        RECT  0.16 -0.28 0.32 0.92 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 3.60 3.48 ;
        RECT  3.14 2.88 3.42 3.48 ;
        RECT  2.56 2.06 2.84 2.66 ;
        RECT  2.62 2.06 2.78 3.48 ;
        RECT  0.10 2.16 0.38 2.44 ;
        RECT  0.16 2.16 0.32 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.64 0.94 0.92 ;
        RECT  0.78 1.46 1.22 1.74 ;
        RECT  0.78 0.64 0.94 2.44 ;
        RECT  0.62 2.16 0.94 2.44 ;
        RECT  1.10 0.64 1.38 0.92 ;
        RECT  2.14 0.64 2.42 0.92 ;
        RECT  1.22 0.64 1.38 1.28 ;
        RECT  2.14 0.64 2.30 1.28 ;
        RECT  1.22 1.12 3.04 1.28 ;
        RECT  2.88 1.12 3.04 1.74 ;
        RECT  2.88 1.46 3.16 1.74 ;
        RECT  1.40 1.12 1.56 2.44 ;
        RECT  1.24 2.16 1.70 2.44 ;
    END
END OR3I1SP2V1_0

MACRO OR3I1SP1V1_0
    CLASS CORE ;
    FOREIGN OR3I1SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.72 1.44 2.04 1.86 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.34 1.46 2.74 1.74 ;
        END
    END IN3
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 6.06  LAYER ME1  ;
        ANTENNADIFFAREA 2.64  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        ANTENNAMAXAREACAR 45.10  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.04 2.16 3.48 2.44 ;
        RECT  3.32 0.64 3.48 2.44 ;
        RECT  3.18 0.64 3.48 0.92 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 3.60 3.48 ;
        RECT  3.14 2.88 3.42 3.48 ;
        RECT  2.52 2.16 2.80 2.44 ;
        RECT  2.58 2.16 2.74 3.48 ;
        RECT  0.10 2.16 0.38 2.44 ;
        RECT  0.16 2.16 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 3.60 0.28 ;
        RECT  3.14 -0.28 3.42 0.32 ;
        RECT  2.66 0.64 2.94 0.92 ;
        RECT  2.72 -0.28 2.88 0.92 ;
        RECT  1.62 0.64 1.90 0.92 ;
        RECT  1.68 -0.28 1.84 0.92 ;
        RECT  0.10 0.64 0.38 0.92 ;
        RECT  0.16 -0.28 0.32 0.92 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.64 0.94 0.92 ;
        RECT  0.78 1.46 1.22 1.74 ;
        RECT  0.78 0.64 0.94 2.44 ;
        RECT  0.62 2.16 0.94 2.44 ;
        RECT  1.10 0.64 1.38 0.92 ;
        RECT  2.14 0.64 2.42 0.92 ;
        RECT  1.22 0.64 1.38 1.28 ;
        RECT  2.14 0.64 2.30 1.28 ;
        RECT  1.22 1.12 3.15 1.28 ;
        RECT  2.87 1.08 3.15 1.36 ;
        RECT  1.40 1.12 1.56 2.44 ;
        RECT  1.24 2.16 1.70 2.44 ;
    END
END OR3I1SP1V1_0

MACRO OR3AND2SP8V1_0
    CLASS CORE ;
    FOREIGN OR3AND2SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 12.04  LAYER ME1  ;
        ANTENNADIFFAREA 6.67  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.71  LAYER ME1  ;
        ANTENNAMAXAREACAR 16.95  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.20 1.97 5.48 2.57 ;
        RECT  5.20 0.63 5.48 1.23 ;
        RECT  5.20 0.63 5.36 2.57 ;
        RECT  4.28 1.52 5.36 1.68 ;
        RECT  4.28 1.46 4.74 1.74 ;
        RECT  4.16 1.97 4.44 2.57 ;
        RECT  4.28 0.63 4.44 2.57 ;
        RECT  4.16 0.63 4.44 1.23 ;
        END
    END OUT
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.32 1.39 3.60 1.81 ;
        END
    END IN4
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.34 1.46 1.94 1.74 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.44 1.14 1.86 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.44 0.38 1.86 ;
        END
    END IN1
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 6.40 0.28 ;
        RECT  5.78 -0.28 6.22 0.32 ;
        RECT  5.72 0.63 6.00 1.23 ;
        RECT  5.78 -0.28 5.94 1.23 ;
        RECT  4.68 0.63 4.96 1.23 ;
        RECT  4.74 -0.28 4.90 1.23 ;
        RECT  3.64 0.63 3.92 0.91 ;
        RECT  3.70 -0.28 3.86 0.91 ;
        RECT  1.66 0.58 1.94 0.86 ;
        RECT  1.72 -0.28 1.88 0.86 ;
        RECT  0.62 0.58 0.90 0.86 ;
        RECT  0.68 -0.28 0.84 0.86 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 6.40 3.48 ;
        RECT  5.78 2.88 6.22 3.48 ;
        RECT  5.72 1.97 6.00 2.57 ;
        RECT  5.78 1.97 5.94 3.48 ;
        RECT  4.68 1.97 4.96 2.57 ;
        RECT  4.74 1.97 4.90 3.48 ;
        RECT  3.64 1.97 3.92 2.57 ;
        RECT  3.70 1.97 3.86 3.48 ;
        RECT  2.56 1.97 2.84 2.25 ;
        RECT  2.62 1.97 2.78 3.48 ;
        RECT  1.52 2.16 1.80 2.44 ;
        RECT  1.58 2.16 1.74 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.58 0.38 0.86 ;
        RECT  1.14 0.58 1.42 0.86 ;
        RECT  0.22 0.58 0.38 1.18 ;
        RECT  1.14 0.58 1.30 1.18 ;
        RECT  0.22 1.02 2.08 1.18 ;
        RECT  1.80 1.02 2.08 1.30 ;
        RECT  0.54 1.02 0.70 2.44 ;
        RECT  0.24 2.16 0.70 2.44 ;
        RECT  2.18 0.58 2.46 0.86 ;
        RECT  2.24 1.46 2.68 1.74 ;
        RECT  2.24 0.58 2.40 2.44 ;
        RECT  2.04 2.16 2.40 2.44 ;
        RECT  2.70 0.63 3.16 0.91 ;
        RECT  3.00 1.07 3.98 1.23 ;
        RECT  3.82 1.07 3.98 1.74 ;
        RECT  3.82 1.46 4.10 1.74 ;
        RECT  3.00 0.63 3.16 2.25 ;
        RECT  3.00 1.97 3.36 2.25 ;
    END
END OR3AND2SP8V1_0

MACRO OR3AND2SP4V1_0
    CLASS CORE ;
    FOREIGN OR3AND2SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 9.71  LAYER ME1  ;
        ANTENNADIFFAREA 4.84  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.42  LAYER ME1  ;
        ANTENNAMAXAREACAR 22.98  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.28 1.46 4.74 1.74 ;
        RECT  4.16 1.97 4.44 2.57 ;
        RECT  4.28 0.63 4.44 2.57 ;
        RECT  4.16 0.63 4.44 1.23 ;
        END
    END OUT
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.32 1.39 3.60 1.81 ;
        END
    END IN4
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.34 1.46 1.94 1.74 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.44 1.14 1.86 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.44 0.38 1.86 ;
        END
    END IN1
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 5.20 0.28 ;
        RECT  4.74 -0.28 5.02 0.32 ;
        RECT  4.68 0.63 4.96 1.23 ;
        RECT  4.74 -0.28 4.90 1.23 ;
        RECT  3.64 0.63 3.92 0.91 ;
        RECT  3.70 -0.28 3.86 0.91 ;
        RECT  1.66 0.58 1.94 0.86 ;
        RECT  1.72 -0.28 1.88 0.86 ;
        RECT  0.62 0.58 0.90 0.86 ;
        RECT  0.68 -0.28 0.84 0.86 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 5.20 3.48 ;
        RECT  4.74 2.88 5.02 3.48 ;
        RECT  4.68 1.97 4.96 2.57 ;
        RECT  4.74 1.97 4.90 3.48 ;
        RECT  3.64 1.97 3.92 2.57 ;
        RECT  3.70 1.97 3.86 3.48 ;
        RECT  2.56 1.97 2.84 2.25 ;
        RECT  2.62 1.97 2.78 3.48 ;
        RECT  1.52 2.16 1.80 2.44 ;
        RECT  1.58 2.16 1.74 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.58 0.38 0.86 ;
        RECT  1.14 0.58 1.42 0.86 ;
        RECT  0.22 0.58 0.38 1.18 ;
        RECT  1.14 0.58 1.30 1.18 ;
        RECT  0.22 1.02 2.08 1.18 ;
        RECT  1.80 1.02 2.08 1.30 ;
        RECT  0.54 1.02 0.70 2.44 ;
        RECT  0.24 2.16 0.70 2.44 ;
        RECT  2.18 0.58 2.46 0.86 ;
        RECT  2.24 1.46 2.68 1.74 ;
        RECT  2.24 0.58 2.40 2.44 ;
        RECT  2.04 2.16 2.40 2.44 ;
        RECT  2.70 0.63 3.16 0.91 ;
        RECT  3.00 1.07 3.98 1.23 ;
        RECT  3.82 1.07 3.98 1.74 ;
        RECT  3.82 1.46 4.10 1.74 ;
        RECT  3.00 0.63 3.16 2.25 ;
        RECT  3.00 1.97 3.36 2.25 ;
    END
END OR3AND2SP4V1_0

MACRO OR3AND2SP2V1_0
    CLASS CORE ;
    FOREIGN OR3AND2SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 8.82  LAYER ME1  ;
        ANTENNADIFFAREA 3.93  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.28  LAYER ME1  ;
        ANTENNAMAXAREACAR 31.67  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.16 1.97 4.68 2.13 ;
        RECT  4.52 1.07 4.68 2.13 ;
        RECT  4.16 1.07 4.68 1.23 ;
        RECT  4.16 1.97 4.44 2.57 ;
        RECT  4.16 0.63 4.44 1.23 ;
        END
    END OUT
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.32 1.39 3.60 1.81 ;
        END
    END IN4
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.34 1.46 1.94 1.74 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.44 1.14 1.86 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.44 0.38 1.86 ;
        END
    END IN1
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.80 0.28 ;
        RECT  4.34 -0.28 4.62 0.32 ;
        RECT  3.64 0.63 3.92 0.91 ;
        RECT  3.70 -0.28 3.86 0.91 ;
        RECT  1.66 0.58 1.94 0.86 ;
        RECT  1.72 -0.28 1.88 0.86 ;
        RECT  0.62 0.58 0.90 0.86 ;
        RECT  0.68 -0.28 0.84 0.86 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.80 3.48 ;
        RECT  4.34 2.88 4.62 3.48 ;
        RECT  3.64 1.97 3.92 2.57 ;
        RECT  3.70 1.97 3.86 3.48 ;
        RECT  2.56 1.97 2.84 2.25 ;
        RECT  2.62 1.97 2.78 3.48 ;
        RECT  1.52 2.16 1.80 2.44 ;
        RECT  1.58 2.16 1.74 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.58 0.38 0.86 ;
        RECT  1.14 0.58 1.42 0.86 ;
        RECT  0.22 0.58 0.38 1.18 ;
        RECT  1.14 0.58 1.30 1.18 ;
        RECT  0.22 1.02 2.08 1.18 ;
        RECT  1.80 1.02 2.08 1.30 ;
        RECT  0.54 1.02 0.70 2.44 ;
        RECT  0.24 2.16 0.70 2.44 ;
        RECT  2.18 0.58 2.46 0.86 ;
        RECT  2.24 1.46 2.68 1.74 ;
        RECT  2.24 0.58 2.40 2.44 ;
        RECT  2.04 2.16 2.40 2.44 ;
        RECT  2.70 0.63 3.16 0.91 ;
        RECT  3.00 1.07 3.98 1.23 ;
        RECT  3.82 1.07 3.98 1.74 ;
        RECT  3.82 1.46 4.10 1.74 ;
        RECT  3.00 0.63 3.16 2.25 ;
        RECT  3.00 1.97 3.36 2.25 ;
    END
END OR3AND2SP2V1_0

MACRO OR3AND2SP1V1_0
    CLASS CORE ;
    FOREIGN OR3AND2SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.44 0.38 1.86 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.44 1.14 1.86 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.34 1.46 1.94 1.74 ;
        END
    END IN3
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 8.18  LAYER ME1  ;
        ANTENNADIFFAREA 3.47  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        ANTENNAMAXAREACAR 40.56  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.12 1.97 4.68 2.13 ;
        RECT  4.52 0.75 4.68 2.13 ;
        RECT  4.12 0.75 4.68 0.91 ;
        RECT  4.12 1.97 4.40 2.25 ;
        RECT  4.12 0.63 4.40 0.91 ;
        END
    END OUT
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.32 1.39 3.60 1.81 ;
        END
    END IN4
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.80 3.48 ;
        RECT  4.34 2.88 4.62 3.48 ;
        RECT  3.60 1.97 3.88 2.25 ;
        RECT  3.66 1.97 3.82 3.48 ;
        RECT  2.56 1.97 2.84 2.25 ;
        RECT  2.62 1.97 2.78 3.48 ;
        RECT  1.52 2.16 1.80 2.44 ;
        RECT  1.58 2.16 1.74 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.80 0.28 ;
        RECT  4.34 -0.28 4.62 0.32 ;
        RECT  3.60 0.63 3.88 0.91 ;
        RECT  3.66 -0.28 3.82 0.91 ;
        RECT  1.66 0.58 1.94 0.86 ;
        RECT  1.72 -0.28 1.88 0.86 ;
        RECT  0.62 0.58 0.90 0.86 ;
        RECT  0.68 -0.28 0.84 0.86 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.58 0.38 0.86 ;
        RECT  1.14 0.58 1.42 0.86 ;
        RECT  0.22 0.58 0.38 1.18 ;
        RECT  1.14 0.58 1.30 1.18 ;
        RECT  0.22 1.02 2.08 1.18 ;
        RECT  1.80 1.02 2.08 1.30 ;
        RECT  0.54 1.02 0.70 2.44 ;
        RECT  0.24 2.16 0.70 2.44 ;
        RECT  2.18 0.58 2.46 0.86 ;
        RECT  2.24 1.46 2.68 1.74 ;
        RECT  2.24 0.58 2.40 2.44 ;
        RECT  2.04 2.16 2.40 2.44 ;
        RECT  2.70 0.63 3.16 0.91 ;
        RECT  3.00 1.08 4.05 1.24 ;
        RECT  3.77 1.07 4.05 1.35 ;
        RECT  3.00 0.63 3.16 2.25 ;
        RECT  3.00 1.97 3.36 2.25 ;
    END
END OR3AND2SP1V1_0

MACRO OR2SP8V1_0
    CLASS CORE ;
    FOREIGN OR2SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 7.06  LAYER ME1  ;
        ANTENNADIFFAREA 4.10  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.58  LAYER ME1  ;
        ANTENNAMAXAREACAR 12.26  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.74 2.02 3.02 2.62 ;
        RECT  1.70 1.04 3.02 1.20 ;
        RECT  2.74 0.92 3.02 1.20 ;
        RECT  1.70 2.02 3.02 2.18 ;
        RECT  2.12 1.04 2.28 2.18 ;
        RECT  1.70 2.02 1.98 2.62 ;
        RECT  1.70 0.92 1.98 1.20 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.00 3.48 ;
        RECT  3.38 2.88 3.82 3.48 ;
        RECT  3.38 2.02 3.54 3.48 ;
        RECT  3.26 2.02 3.54 2.62 ;
        RECT  2.22 2.34 2.50 2.62 ;
        RECT  2.28 2.34 2.44 3.48 ;
        RECT  1.18 2.02 1.46 2.62 ;
        RECT  1.24 2.02 1.40 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.00 0.28 ;
        RECT  3.38 -0.28 3.82 0.32 ;
        RECT  3.26 0.60 3.54 0.88 ;
        RECT  3.38 -0.28 3.54 0.88 ;
        RECT  2.22 0.60 2.50 0.88 ;
        RECT  2.28 -0.28 2.44 0.88 ;
        RECT  1.18 0.60 1.46 0.88 ;
        RECT  1.24 -0.28 1.40 0.88 ;
        RECT  0.10 0.63 0.38 0.91 ;
        RECT  0.16 -0.28 0.32 0.91 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.54 0.63 0.90 0.91 ;
        RECT  0.54 1.07 1.50 1.23 ;
        RECT  1.34 1.07 1.50 1.62 ;
        RECT  1.34 1.34 1.62 1.62 ;
        RECT  0.54 0.63 0.70 2.18 ;
        RECT  0.24 2.02 0.70 2.18 ;
        RECT  0.24 2.02 0.52 2.30 ;
    END
END OR2SP8V1_0

MACRO OR2SP4V1_0
    CLASS CORE ;
    FOREIGN OR2SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 2.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 4.59  LAYER ME1  ;
        ANTENNADIFFAREA 2.76  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.29  LAYER ME1  ;
        ANTENNAMAXAREACAR 15.92  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.82 1.52 2.28 1.68 ;
        RECT  1.70 2.02 1.98 2.62 ;
        RECT  1.82 0.92 1.98 2.62 ;
        RECT  1.70 0.92 1.98 1.20 ;
        END
    END OUT
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 2.80 3.48 ;
        RECT  2.28 2.88 2.62 3.48 ;
        RECT  2.22 2.02 2.50 2.62 ;
        RECT  2.28 2.02 2.44 3.48 ;
        RECT  1.18 2.02 1.46 2.62 ;
        RECT  1.24 2.02 1.40 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 2.80 0.28 ;
        RECT  2.28 -0.28 2.62 0.32 ;
        RECT  2.22 0.60 2.50 0.88 ;
        RECT  2.28 -0.28 2.44 0.88 ;
        RECT  1.18 0.60 1.46 0.88 ;
        RECT  1.24 -0.28 1.40 0.88 ;
        RECT  0.10 0.63 0.38 0.91 ;
        RECT  0.16 -0.28 0.32 0.91 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.54 0.63 0.90 0.91 ;
        RECT  0.54 1.07 1.50 1.23 ;
        RECT  1.34 1.07 1.50 1.62 ;
        RECT  1.34 1.34 1.62 1.62 ;
        RECT  0.54 0.63 0.70 2.18 ;
        RECT  0.24 2.02 0.70 2.18 ;
        RECT  0.24 2.02 0.52 2.30 ;
    END
END OR2SP4V1_0

MACRO OR2SP2V1_0
    CLASS CORE ;
    FOREIGN OR2SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 2.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 3.80  LAYER ME1  ;
        ANTENNADIFFAREA 2.15  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.14  LAYER ME1  ;
        ANTENNAMAXAREACAR 26.39  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.70 2.02 2.28 2.18 ;
        RECT  2.12 1.04 2.28 2.18 ;
        RECT  1.70 1.04 2.28 1.20 ;
        RECT  1.70 2.02 1.98 2.62 ;
        RECT  1.70 0.92 1.98 1.20 ;
        END
    END OUT
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 2.40 0.28 ;
        RECT  1.94 -0.28 2.22 0.32 ;
        RECT  1.18 0.60 1.46 0.88 ;
        RECT  1.24 -0.28 1.40 0.88 ;
        RECT  0.10 0.63 0.38 0.91 ;
        RECT  0.16 -0.28 0.32 0.91 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 2.40 3.48 ;
        RECT  1.94 2.88 2.22 3.48 ;
        RECT  1.18 2.02 1.46 2.62 ;
        RECT  1.24 2.02 1.40 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.54 0.63 0.90 0.91 ;
        RECT  0.54 1.07 1.50 1.23 ;
        RECT  1.34 1.07 1.50 1.62 ;
        RECT  1.34 1.34 1.62 1.62 ;
        RECT  0.54 0.63 0.70 2.18 ;
        RECT  0.24 2.02 0.70 2.18 ;
        RECT  0.24 2.02 0.52 2.30 ;
    END
END OR2SP2V1_0

MACRO OR2SP1V1_0
    CLASS CORE ;
    FOREIGN OR2SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 2.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 3.73  LAYER ME1  ;
        ANTENNADIFFAREA 1.69  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 55.57  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.66 0.63 1.94 0.91 ;
        RECT  1.57 2.02 1.92 2.30 ;
        RECT  1.76 0.63 1.92 2.30 ;
        RECT  1.72 1.52 1.92 1.68 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 2.40 3.48 ;
        RECT  1.94 2.88 2.22 3.48 ;
        RECT  1.05 2.02 1.33 2.30 ;
        RECT  1.11 2.02 1.27 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 2.40 0.28 ;
        RECT  1.94 -0.28 2.22 0.32 ;
        RECT  1.14 0.63 1.42 0.91 ;
        RECT  1.20 -0.28 1.36 0.91 ;
        RECT  0.10 0.63 0.38 0.91 ;
        RECT  0.16 -0.28 0.32 0.91 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.54 0.63 0.90 0.91 ;
        RECT  0.54 1.07 1.60 1.23 ;
        RECT  1.32 1.07 1.60 1.35 ;
        RECT  0.54 0.63 0.70 2.18 ;
        RECT  0.15 2.02 0.70 2.18 ;
        RECT  0.15 2.02 0.43 2.30 ;
    END
END OR2SP1V1_0

MACRO OR2NAND3SP8V1_0
    CLASS CORE ;
    FOREIGN OR2NAND3SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.39 0.70 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.16 1.81 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.32 1.39 1.64 1.81 ;
        END
    END IN3
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 14.14  LAYER ME1  ;
        ANTENNADIFFAREA 7.27  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.78  LAYER ME1  ;
        ANTENNAMAXAREACAR 18.18  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.38 1.90 6.66 2.50 ;
        RECT  6.38 0.64 6.66 1.24 ;
        RECT  6.38 0.64 6.54 2.50 ;
        RECT  5.26 1.52 6.54 1.68 ;
        RECT  5.32 1.90 5.62 2.50 ;
        RECT  5.32 0.64 5.62 1.24 ;
        RECT  5.26 1.46 5.54 1.74 ;
        RECT  5.32 0.64 5.48 2.50 ;
        END
    END OUT
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.12 1.44 2.40 1.83 ;
        END
    END IN4
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 7.60 0.28 ;
        RECT  6.98 -0.28 7.42 0.32 ;
        RECT  6.90 0.64 7.18 1.24 ;
        RECT  6.98 -0.28 7.14 1.24 ;
        RECT  5.86 0.64 6.14 1.24 ;
        RECT  5.92 -0.28 6.08 1.24 ;
        RECT  4.82 0.64 5.10 1.24 ;
        RECT  4.88 -0.28 5.04 1.24 ;
        RECT  3.82 0.68 4.10 0.96 ;
        RECT  3.88 -0.28 4.04 0.96 ;
        RECT  2.78 0.68 3.06 0.96 ;
        RECT  2.84 -0.28 3.00 0.96 ;
        RECT  1.14 0.60 1.42 0.88 ;
        RECT  1.20 -0.28 1.36 0.88 ;
        RECT  0.10 0.60 0.38 0.88 ;
        RECT  0.16 -0.28 0.32 0.88 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 7.60 3.48 ;
        RECT  6.98 2.88 7.42 3.48 ;
        RECT  6.90 1.90 7.18 2.50 ;
        RECT  6.98 1.90 7.14 3.48 ;
        RECT  5.86 1.90 6.14 2.50 ;
        RECT  5.92 1.90 6.08 3.48 ;
        RECT  4.82 1.90 5.10 2.50 ;
        RECT  4.88 1.90 5.04 3.48 ;
        RECT  2.88 2.02 3.16 2.30 ;
        RECT  2.94 2.02 3.10 3.48 ;
        RECT  1.14 2.02 1.42 2.30 ;
        RECT  1.20 2.02 1.36 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.60 0.90 0.88 ;
        RECT  0.62 0.60 0.78 1.23 ;
        RECT  0.08 1.07 0.78 1.23 ;
        RECT  0.08 2.02 0.52 2.30 ;
        RECT  0.08 1.07 0.24 2.76 ;
        RECT  0.08 2.48 0.38 2.76 ;
        RECT  1.66 0.60 1.96 0.88 ;
        RECT  1.80 0.98 2.08 1.26 ;
        RECT  1.80 0.60 1.96 2.30 ;
        RECT  1.66 2.02 1.96 2.30 ;
        RECT  2.26 0.68 2.54 0.96 ;
        RECT  2.38 0.68 2.54 1.28 ;
        RECT  2.38 1.12 3.20 1.28 ;
        RECT  3.04 1.12 3.20 1.71 ;
        RECT  3.04 1.43 3.32 1.71 ;
        RECT  2.56 1.12 2.72 2.30 ;
        RECT  2.36 2.02 2.72 2.30 ;
        RECT  3.30 0.68 3.58 0.96 ;
        RECT  4.34 0.68 4.62 0.96 ;
        RECT  3.42 0.68 3.58 1.28 ;
        RECT  3.42 1.12 4.50 1.28 ;
        RECT  4.34 1.52 5.10 1.68 ;
        RECT  4.82 1.46 5.10 1.74 ;
        RECT  4.34 0.68 4.50 2.30 ;
        RECT  4.16 2.02 4.50 2.30 ;
    END
END OR2NAND3SP8V1_0

MACRO OR2NAND3SP4V1_0
    CLASS CORE ;
    FOREIGN OR2NAND3SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.12 1.44 2.40 1.83 ;
        END
    END IN4
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 11.75  LAYER ME1  ;
        ANTENNADIFFAREA 5.45  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER ME1  ;
        ANTENNAMAXAREACAR 23.99  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.32 1.90 5.62 2.50 ;
        RECT  5.32 0.64 5.62 1.24 ;
        RECT  5.26 1.46 5.54 1.74 ;
        RECT  5.32 0.64 5.48 2.50 ;
        END
    END OUT
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.32 1.39 1.64 1.81 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.16 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.39 0.70 1.81 ;
        END
    END IN1
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 6.40 0.28 ;
        RECT  5.92 -0.28 6.22 0.32 ;
        RECT  5.86 0.64 6.14 1.24 ;
        RECT  5.92 -0.28 6.08 1.24 ;
        RECT  4.82 0.64 5.10 1.24 ;
        RECT  4.88 -0.28 5.04 1.24 ;
        RECT  3.82 0.68 4.10 0.96 ;
        RECT  3.88 -0.28 4.04 0.96 ;
        RECT  2.78 0.68 3.06 0.96 ;
        RECT  2.84 -0.28 3.00 0.96 ;
        RECT  1.14 0.60 1.42 0.88 ;
        RECT  1.20 -0.28 1.36 0.88 ;
        RECT  0.10 0.60 0.38 0.88 ;
        RECT  0.16 -0.28 0.32 0.88 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 6.40 3.48 ;
        RECT  5.92 2.88 6.22 3.48 ;
        RECT  5.86 1.90 6.14 2.50 ;
        RECT  5.92 1.90 6.08 3.48 ;
        RECT  4.82 1.90 5.10 2.50 ;
        RECT  4.88 1.90 5.04 3.48 ;
        RECT  2.88 2.02 3.16 2.30 ;
        RECT  2.94 2.02 3.10 3.48 ;
        RECT  1.14 2.02 1.42 2.30 ;
        RECT  1.20 2.02 1.36 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.60 0.90 0.88 ;
        RECT  0.62 0.60 0.78 1.23 ;
        RECT  0.08 1.07 0.78 1.23 ;
        RECT  0.08 2.02 0.52 2.30 ;
        RECT  0.08 1.07 0.24 2.76 ;
        RECT  0.08 2.48 0.38 2.76 ;
        RECT  1.66 0.60 1.96 0.88 ;
        RECT  1.80 0.98 2.08 1.26 ;
        RECT  1.80 0.60 1.96 2.30 ;
        RECT  1.66 2.02 1.96 2.30 ;
        RECT  2.26 0.68 2.54 0.96 ;
        RECT  2.38 0.68 2.54 1.28 ;
        RECT  2.38 1.12 3.20 1.28 ;
        RECT  3.04 1.12 3.20 1.71 ;
        RECT  3.04 1.43 3.32 1.71 ;
        RECT  2.56 1.12 2.72 2.30 ;
        RECT  2.36 2.02 2.72 2.30 ;
        RECT  3.30 0.68 3.58 0.96 ;
        RECT  4.34 0.68 4.62 0.96 ;
        RECT  3.42 0.68 3.58 1.28 ;
        RECT  3.42 1.12 4.50 1.28 ;
        RECT  4.34 1.52 5.10 1.68 ;
        RECT  4.82 1.46 5.10 1.74 ;
        RECT  4.34 0.68 4.50 2.30 ;
        RECT  4.16 2.02 4.50 2.30 ;
    END
END OR2NAND3SP4V1_0

MACRO OR2NAND3SP2V1_0
    CLASS CORE ;
    FOREIGN OR2NAND3SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 10.84  LAYER ME1  ;
        ANTENNADIFFAREA 4.84  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.35  LAYER ME1  ;
        ANTENNAMAXAREACAR 31.35  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.32 1.90 5.62 2.50 ;
        RECT  5.32 0.64 5.62 1.24 ;
        RECT  5.26 1.46 5.54 1.74 ;
        RECT  5.32 0.64 5.48 2.50 ;
        END
    END OUT
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.12 1.71 2.40 2.08 ;
        END
    END IN4
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.32 1.39 1.64 1.81 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.16 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.39 0.70 1.81 ;
        END
    END IN1
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 6.00 3.48 ;
        RECT  5.54 2.88 5.82 3.48 ;
        RECT  4.82 1.90 5.10 2.50 ;
        RECT  4.88 1.90 5.04 3.48 ;
        RECT  2.88 2.24 3.16 2.52 ;
        RECT  2.94 2.24 3.10 3.48 ;
        RECT  1.14 2.02 1.42 2.30 ;
        RECT  1.20 2.02 1.36 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 6.00 0.28 ;
        RECT  5.54 -0.28 5.82 0.32 ;
        RECT  4.82 0.64 5.10 1.24 ;
        RECT  4.88 -0.28 5.04 1.24 ;
        RECT  3.82 0.68 4.10 0.96 ;
        RECT  3.88 -0.28 4.04 0.96 ;
        RECT  2.78 0.68 3.06 0.96 ;
        RECT  2.84 -0.28 3.00 0.96 ;
        RECT  1.14 0.63 1.42 0.91 ;
        RECT  1.20 -0.28 1.36 0.91 ;
        RECT  0.10 0.63 0.38 0.91 ;
        RECT  0.16 -0.28 0.32 0.91 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.63 0.90 0.91 ;
        RECT  0.62 0.63 0.78 1.23 ;
        RECT  0.08 1.07 0.78 1.23 ;
        RECT  0.08 2.02 0.52 2.30 ;
        RECT  0.08 1.07 0.24 2.76 ;
        RECT  0.08 2.48 0.38 2.76 ;
        RECT  1.66 0.63 1.96 0.91 ;
        RECT  1.80 1.01 2.08 1.29 ;
        RECT  1.80 0.63 1.96 2.30 ;
        RECT  1.66 2.02 1.96 2.30 ;
        RECT  2.26 0.68 2.54 0.96 ;
        RECT  2.38 0.68 2.54 1.28 ;
        RECT  2.38 1.12 2.72 1.28 ;
        RECT  2.56 1.49 3.32 1.65 ;
        RECT  3.04 1.43 3.32 1.71 ;
        RECT  2.56 1.12 2.72 2.52 ;
        RECT  2.36 2.24 2.72 2.52 ;
        RECT  3.30 0.68 3.58 0.96 ;
        RECT  4.34 0.68 4.62 0.96 ;
        RECT  3.42 0.68 3.58 1.28 ;
        RECT  3.42 1.12 4.50 1.28 ;
        RECT  4.34 1.52 5.10 1.68 ;
        RECT  4.82 1.46 5.10 1.74 ;
        RECT  4.34 0.68 4.50 2.52 ;
        RECT  4.16 2.24 4.50 2.52 ;
    END
END OR2NAND3SP2V1_0

MACRO OR2NAND3SP1V1_0
    CLASS CORE ;
    FOREIGN OR2NAND3SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.39 0.70 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.16 1.81 ;
        END
    END IN2
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.12 1.44 2.40 1.83 ;
        END
    END IN4
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 10.27  LAYER ME1  ;
        ANTENNADIFFAREA 4.41  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.27  LAYER ME1  ;
        ANTENNAMAXAREACAR 38.22  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.32 1.90 5.62 2.18 ;
        RECT  5.32 0.96 5.62 1.24 ;
        RECT  5.26 1.46 5.54 1.74 ;
        RECT  5.32 0.96 5.48 2.18 ;
        END
    END OUT
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.32 1.39 1.64 1.81 ;
        END
    END IN3
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 6.00 3.48 ;
        RECT  5.54 2.88 5.82 3.48 ;
        RECT  4.82 1.90 5.10 2.18 ;
        RECT  4.88 1.90 5.04 3.48 ;
        RECT  2.88 2.02 3.16 2.30 ;
        RECT  2.94 2.02 3.10 3.48 ;
        RECT  1.14 2.02 1.42 2.30 ;
        RECT  1.20 2.02 1.36 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 6.00 0.28 ;
        RECT  5.54 -0.28 5.82 0.32 ;
        RECT  4.82 0.96 5.10 1.24 ;
        RECT  4.88 -0.28 5.04 1.24 ;
        RECT  3.82 0.68 4.10 0.96 ;
        RECT  3.88 -0.28 4.04 0.96 ;
        RECT  2.78 0.68 3.06 0.96 ;
        RECT  2.84 -0.28 3.00 0.96 ;
        RECT  1.14 0.60 1.42 0.88 ;
        RECT  1.20 -0.28 1.36 0.88 ;
        RECT  0.10 0.60 0.38 0.88 ;
        RECT  0.16 -0.28 0.32 0.88 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.60 0.90 0.88 ;
        RECT  0.62 0.60 0.78 1.23 ;
        RECT  0.08 1.07 0.78 1.23 ;
        RECT  0.08 2.02 0.52 2.30 ;
        RECT  0.08 1.07 0.24 2.76 ;
        RECT  0.08 2.48 0.38 2.76 ;
        RECT  1.66 0.60 1.96 0.88 ;
        RECT  1.80 0.98 2.08 1.26 ;
        RECT  1.80 0.60 1.96 2.30 ;
        RECT  1.66 2.02 1.96 2.30 ;
        RECT  2.26 0.68 2.54 0.96 ;
        RECT  2.38 0.68 2.54 1.28 ;
        RECT  2.38 1.12 3.20 1.28 ;
        RECT  3.04 1.12 3.20 1.71 ;
        RECT  3.04 1.43 3.32 1.71 ;
        RECT  2.56 1.12 2.72 2.30 ;
        RECT  2.36 2.02 2.72 2.30 ;
        RECT  3.30 0.68 3.58 0.96 ;
        RECT  4.34 0.68 4.62 0.96 ;
        RECT  3.42 0.68 3.58 1.28 ;
        RECT  3.42 1.12 4.50 1.28 ;
        RECT  4.34 1.52 5.10 1.68 ;
        RECT  4.82 1.46 5.10 1.74 ;
        RECT  4.34 0.68 4.50 2.30 ;
        RECT  4.16 2.02 4.50 2.30 ;
    END
END OR2NAND3SP1V1_0

MACRO OR2NAND2SP8V1_0
    CLASS CORE ;
    FOREIGN OR2NAND2SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 11.33  LAYER ME1  ;
        ANTENNADIFFAREA 6.34  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.71  LAYER ME1  ;
        ANTENNAMAXAREACAR 15.95  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.83 1.98 5.11 2.58 ;
        RECT  4.83 0.64 5.11 1.24 ;
        RECT  4.83 0.64 4.99 2.58 ;
        RECT  3.87 1.52 4.99 1.68 ;
        RECT  3.87 1.46 4.34 1.74 ;
        RECT  3.79 1.98 4.07 2.58 ;
        RECT  3.79 0.64 4.07 1.24 ;
        RECT  3.87 0.64 4.03 2.58 ;
        END
    END OUT
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.32 1.39 1.64 1.81 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.16 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.39 0.70 1.81 ;
        END
    END IN1
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 6.00 0.28 ;
        RECT  5.41 -0.28 5.82 0.32 ;
        RECT  5.35 0.64 5.63 1.24 ;
        RECT  5.41 -0.28 5.57 1.24 ;
        RECT  4.31 0.64 4.59 1.24 ;
        RECT  4.37 -0.28 4.53 1.24 ;
        RECT  3.27 0.64 3.55 1.24 ;
        RECT  3.33 -0.28 3.49 1.24 ;
        RECT  2.19 0.96 2.47 1.24 ;
        RECT  2.25 -0.28 2.41 1.24 ;
        RECT  1.19 0.63 1.47 0.91 ;
        RECT  1.25 -0.28 1.41 0.91 ;
        RECT  0.15 0.63 0.43 0.91 ;
        RECT  0.21 -0.28 0.37 0.91 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 6.00 3.48 ;
        RECT  5.41 2.88 5.82 3.48 ;
        RECT  5.35 1.98 5.63 2.58 ;
        RECT  5.41 1.98 5.57 3.48 ;
        RECT  4.31 1.98 4.59 2.58 ;
        RECT  4.37 1.98 4.53 3.48 ;
        RECT  3.27 1.98 3.55 2.58 ;
        RECT  3.33 1.98 3.49 3.48 ;
        RECT  1.14 2.02 1.42 2.30 ;
        RECT  1.20 2.02 1.36 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.67 0.63 0.95 0.91 ;
        RECT  0.67 0.63 0.83 1.23 ;
        RECT  0.08 1.07 0.83 1.23 ;
        RECT  0.08 2.02 0.52 2.30 ;
        RECT  0.08 1.07 0.24 2.76 ;
        RECT  0.08 2.48 0.38 2.76 ;
        RECT  1.71 0.63 1.99 0.91 ;
        RECT  1.80 1.52 2.53 1.68 ;
        RECT  2.25 1.46 2.53 1.74 ;
        RECT  1.80 0.63 1.96 2.30 ;
        RECT  1.66 2.02 1.96 2.30 ;
        RECT  2.71 0.96 2.99 1.24 ;
        RECT  2.77 1.52 3.69 1.68 ;
        RECT  3.41 1.46 3.69 1.74 ;
        RECT  2.77 0.96 2.93 2.18 ;
        RECT  2.33 2.02 2.93 2.18 ;
        RECT  2.33 2.02 2.61 2.30 ;
    END
END OR2NAND2SP8V1_0

MACRO OR2NAND2SP4V1_0
    CLASS CORE ;
    FOREIGN OR2NAND2SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.39 0.70 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.16 1.81 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.32 1.39 1.64 1.81 ;
        END
    END IN3
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 9.00  LAYER ME1  ;
        ANTENNADIFFAREA 4.51  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.42  LAYER ME1  ;
        ANTENNAMAXAREACAR 21.30  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.87 1.46 4.34 1.74 ;
        RECT  3.79 1.98 4.07 2.58 ;
        RECT  3.79 0.64 4.07 1.24 ;
        RECT  3.87 0.64 4.03 2.58 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.80 3.48 ;
        RECT  4.34 2.88 4.62 3.48 ;
        RECT  4.31 1.98 4.59 2.58 ;
        RECT  4.37 1.98 4.53 3.48 ;
        RECT  3.27 1.98 3.55 2.58 ;
        RECT  3.33 1.98 3.49 3.48 ;
        RECT  1.14 2.02 1.42 2.30 ;
        RECT  1.20 2.02 1.36 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.80 0.28 ;
        RECT  4.34 -0.28 4.62 0.32 ;
        RECT  4.31 0.64 4.59 1.24 ;
        RECT  4.37 -0.28 4.53 1.24 ;
        RECT  3.27 0.64 3.55 1.24 ;
        RECT  3.33 -0.28 3.49 1.24 ;
        RECT  2.19 0.96 2.47 1.24 ;
        RECT  2.25 -0.28 2.41 1.24 ;
        RECT  1.19 0.63 1.47 0.91 ;
        RECT  1.25 -0.28 1.41 0.91 ;
        RECT  0.15 0.63 0.43 0.91 ;
        RECT  0.21 -0.28 0.37 0.91 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.67 0.63 0.95 0.91 ;
        RECT  0.67 0.63 0.83 1.23 ;
        RECT  0.08 1.07 0.83 1.23 ;
        RECT  0.08 2.02 0.52 2.30 ;
        RECT  0.08 1.07 0.24 2.76 ;
        RECT  0.08 2.48 0.38 2.76 ;
        RECT  1.71 0.63 1.99 0.91 ;
        RECT  1.80 1.52 2.53 1.68 ;
        RECT  2.25 1.46 2.53 1.74 ;
        RECT  1.80 0.63 1.96 2.30 ;
        RECT  1.66 2.02 1.96 2.30 ;
        RECT  2.71 0.96 2.99 1.24 ;
        RECT  2.77 1.52 3.69 1.68 ;
        RECT  3.41 1.46 3.69 1.74 ;
        RECT  2.77 0.96 2.93 2.18 ;
        RECT  2.33 2.02 2.93 2.18 ;
        RECT  2.33 2.02 2.61 2.30 ;
    END
END OR2NAND2SP4V1_0

MACRO OR2NAND2SP2V1_0
    CLASS CORE ;
    FOREIGN OR2NAND2SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 8.11  LAYER ME1  ;
        ANTENNADIFFAREA 3.69  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.28  LAYER ME1  ;
        ANTENNAMAXAREACAR 29.12  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.87 1.46 4.32 1.74 ;
        RECT  3.79 1.98 4.07 2.58 ;
        RECT  3.79 0.64 4.07 1.24 ;
        RECT  3.87 0.64 4.03 2.58 ;
        END
    END OUT
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.32 1.39 1.64 1.81 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.16 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.39 0.70 1.81 ;
        END
    END IN1
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.40 0.28 ;
        RECT  3.94 -0.28 4.22 0.32 ;
        RECT  3.27 0.64 3.55 1.24 ;
        RECT  3.33 -0.28 3.49 1.24 ;
        RECT  2.19 0.96 2.47 1.24 ;
        RECT  2.25 -0.28 2.41 1.24 ;
        RECT  1.19 0.63 1.47 0.91 ;
        RECT  1.25 -0.28 1.41 0.91 ;
        RECT  0.15 0.63 0.43 0.91 ;
        RECT  0.21 -0.28 0.37 0.91 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.40 3.48 ;
        RECT  3.94 2.88 4.22 3.48 ;
        RECT  3.27 1.98 3.55 2.58 ;
        RECT  3.33 1.98 3.49 3.48 ;
        RECT  1.14 2.02 1.42 2.30 ;
        RECT  1.20 2.02 1.36 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.67 0.63 0.95 0.91 ;
        RECT  0.67 0.63 0.83 1.23 ;
        RECT  0.08 1.07 0.83 1.23 ;
        RECT  0.08 2.02 0.52 2.30 ;
        RECT  0.08 1.07 0.24 2.76 ;
        RECT  0.08 2.48 0.38 2.76 ;
        RECT  1.71 0.63 1.99 0.91 ;
        RECT  1.80 1.52 2.53 1.68 ;
        RECT  2.25 1.46 2.53 1.74 ;
        RECT  1.80 0.63 1.96 2.30 ;
        RECT  1.66 2.02 1.96 2.30 ;
        RECT  2.71 0.96 2.99 1.24 ;
        RECT  2.77 1.52 3.69 1.68 ;
        RECT  3.41 1.46 3.69 1.74 ;
        RECT  2.77 0.96 2.93 2.18 ;
        RECT  2.33 2.02 2.93 2.18 ;
        RECT  2.33 2.02 2.61 2.30 ;
    END
END OR2NAND2SP2V1_0

MACRO OR2NAND2SP1V1_0
    CLASS CORE ;
    FOREIGN OR2NAND2SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.39 0.70 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.16 1.81 ;
        END
    END IN2
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 7.49  LAYER ME1  ;
        ANTENNADIFFAREA 3.23  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        ANTENNAMAXAREACAR 37.14  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.87 1.46 4.32 1.74 ;
        RECT  3.75 2.02 4.03 2.30 ;
        RECT  3.87 0.96 4.03 2.30 ;
        RECT  3.75 0.96 4.03 1.24 ;
        END
    END OUT
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.32 1.39 1.64 1.81 ;
        END
    END IN3
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.40 3.48 ;
        RECT  3.94 2.88 4.22 3.48 ;
        RECT  3.23 2.02 3.51 2.30 ;
        RECT  3.29 2.02 3.45 3.48 ;
        RECT  1.14 2.02 1.42 2.30 ;
        RECT  1.20 2.02 1.36 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.40 0.28 ;
        RECT  3.94 -0.28 4.22 0.32 ;
        RECT  3.23 0.96 3.51 1.24 ;
        RECT  3.29 -0.28 3.45 1.24 ;
        RECT  2.19 0.96 2.47 1.24 ;
        RECT  2.25 -0.28 2.41 1.24 ;
        RECT  1.19 0.63 1.47 0.91 ;
        RECT  1.25 -0.28 1.41 0.91 ;
        RECT  0.15 0.63 0.43 0.91 ;
        RECT  0.21 -0.28 0.37 0.91 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.67 0.63 0.95 0.91 ;
        RECT  0.67 0.63 0.83 1.23 ;
        RECT  0.08 1.07 0.83 1.23 ;
        RECT  0.08 2.02 0.52 2.30 ;
        RECT  0.08 1.07 0.24 2.76 ;
        RECT  0.08 2.48 0.38 2.76 ;
        RECT  1.71 0.63 1.99 0.91 ;
        RECT  1.80 1.52 2.53 1.68 ;
        RECT  2.25 1.46 2.53 1.74 ;
        RECT  1.80 0.63 1.96 2.30 ;
        RECT  1.66 2.02 1.96 2.30 ;
        RECT  2.71 0.96 2.99 1.24 ;
        RECT  2.77 1.52 3.69 1.68 ;
        RECT  3.41 1.46 3.69 1.74 ;
        RECT  2.77 0.96 2.93 2.18 ;
        RECT  2.33 2.02 2.93 2.18 ;
        RECT  2.33 2.02 2.61 2.30 ;
    END
END OR2NAND2SP1V1_0

MACRO OR2I1SP8V1_0
    CLASS CORE ;
    FOREIGN OR2I1SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 8.53  LAYER ME1  ;
        ANTENNADIFFAREA 4.53  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.64  LAYER ME1  ;
        ANTENNAMAXAREACAR 13.27  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.46 1.04 3.78 1.20 ;
        RECT  3.50 0.60 3.78 1.20 ;
        RECT  3.41 2.00 3.69 2.60 ;
        RECT  2.37 2.00 3.69 2.16 ;
        RECT  2.46 0.60 2.74 1.20 ;
        RECT  2.37 2.00 2.68 2.60 ;
        RECT  2.52 0.60 2.68 2.60 ;
        END
    END OUT
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.60 1.45 1.88 1.84 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.43 1.79 0.71 2.21 ;
        END
    END IN1
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.40 0.28 ;
        RECT  4.02 0.60 4.30 1.20 ;
        RECT  4.08 -0.28 4.24 1.20 ;
        RECT  3.94 -0.28 4.24 0.32 ;
        RECT  2.98 0.60 3.26 0.88 ;
        RECT  3.04 -0.28 3.20 0.88 ;
        RECT  1.94 0.60 2.22 0.88 ;
        RECT  2.00 -0.28 2.16 0.88 ;
        RECT  0.86 0.63 1.14 0.91 ;
        RECT  0.92 -0.28 1.08 0.91 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.40 3.48 ;
        RECT  3.94 2.88 4.22 3.48 ;
        RECT  3.93 2.00 4.21 2.60 ;
        RECT  4.02 2.00 4.18 3.48 ;
        RECT  2.89 2.32 3.17 2.60 ;
        RECT  2.98 2.32 3.14 3.48 ;
        RECT  1.85 2.00 2.13 2.60 ;
        RECT  1.91 2.00 2.07 3.48 ;
        RECT  0.62 2.48 0.90 2.76 ;
        RECT  0.68 2.48 0.84 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.34 0.63 0.62 0.91 ;
        RECT  0.11 0.75 0.62 0.91 ;
        RECT  0.11 1.07 1.00 1.23 ;
        RECT  0.84 1.07 1.00 1.63 ;
        RECT  0.84 1.35 1.12 1.63 ;
        RECT  0.11 0.75 0.27 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  1.38 0.63 1.66 0.91 ;
        RECT  1.44 0.63 1.60 1.23 ;
        RECT  1.28 1.07 2.24 1.23 ;
        RECT  2.08 1.07 2.24 1.61 ;
        RECT  2.08 1.33 2.36 1.61 ;
        RECT  1.28 1.07 1.44 2.16 ;
        RECT  0.91 2.00 1.44 2.16 ;
        RECT  0.91 2.00 1.19 2.28 ;
    END
END OR2I1SP8V1_0

MACRO OR2I1SP4V1_0
    CLASS CORE ;
    FOREIGN OR2I1SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.43 1.79 0.71 2.21 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.60 1.45 1.88 1.84 ;
        END
    END IN2
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 6.33  LAYER ME1  ;
        ANTENNADIFFAREA 3.32  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.36  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.82  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.46 0.60 2.74 1.20 ;
        RECT  2.37 2.00 2.68 2.60 ;
        RECT  2.52 0.60 2.68 2.60 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 3.60 3.48 ;
        RECT  2.98 2.88 3.42 3.48 ;
        RECT  2.89 2.00 3.17 2.60 ;
        RECT  2.98 2.00 3.14 3.48 ;
        RECT  1.85 2.00 2.13 2.60 ;
        RECT  1.91 2.00 2.07 3.48 ;
        RECT  0.62 2.48 0.90 2.76 ;
        RECT  0.68 2.48 0.84 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 3.60 0.28 ;
        RECT  3.04 -0.28 3.42 0.32 ;
        RECT  2.98 0.60 3.26 1.20 ;
        RECT  3.04 -0.28 3.20 1.20 ;
        RECT  1.94 0.60 2.22 0.88 ;
        RECT  2.00 -0.28 2.16 0.88 ;
        RECT  0.86 0.63 1.14 0.91 ;
        RECT  0.92 -0.28 1.08 0.91 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.34 0.63 0.62 0.91 ;
        RECT  0.11 0.75 0.62 0.91 ;
        RECT  0.11 1.07 1.00 1.23 ;
        RECT  0.84 1.07 1.00 1.63 ;
        RECT  0.84 1.35 1.12 1.63 ;
        RECT  0.11 0.75 0.27 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  1.38 0.63 1.66 0.91 ;
        RECT  1.44 0.63 1.60 1.23 ;
        RECT  1.28 1.07 2.24 1.23 ;
        RECT  2.08 1.07 2.24 1.61 ;
        RECT  2.08 1.33 2.36 1.61 ;
        RECT  1.28 1.07 1.44 2.16 ;
        RECT  0.91 2.00 1.44 2.16 ;
        RECT  0.91 2.00 1.19 2.28 ;
    END
END OR2I1SP4V1_0

MACRO OR2I1SP2V1_0
    CLASS CORE ;
    FOREIGN OR2I1SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 2.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 5.00  LAYER ME1  ;
        ANTENNADIFFAREA 2.58  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.21  LAYER ME1  ;
        ANTENNAMAXAREACAR 23.67  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.46 0.60 2.74 1.20 ;
        RECT  2.37 2.00 2.68 2.60 ;
        RECT  2.52 0.60 2.68 2.60 ;
        END
    END OUT
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.60 1.45 1.88 1.84 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.43 1.79 0.71 2.21 ;
        END
    END IN1
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 2.80 0.28 ;
        RECT  2.34 -0.28 2.62 0.32 ;
        RECT  1.94 0.60 2.22 0.88 ;
        RECT  2.00 -0.28 2.16 0.88 ;
        RECT  0.86 0.63 1.14 0.91 ;
        RECT  0.92 -0.28 1.08 0.91 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 2.80 3.48 ;
        RECT  2.34 2.88 2.62 3.48 ;
        RECT  1.85 2.00 2.13 2.60 ;
        RECT  1.91 2.00 2.07 3.48 ;
        RECT  0.62 2.48 0.90 2.76 ;
        RECT  0.68 2.48 0.84 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.34 0.63 0.62 0.91 ;
        RECT  0.11 0.75 0.62 0.91 ;
        RECT  0.11 1.07 1.00 1.23 ;
        RECT  0.84 1.07 1.00 1.63 ;
        RECT  0.84 1.35 1.12 1.63 ;
        RECT  0.11 0.75 0.27 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  1.38 0.63 1.66 0.91 ;
        RECT  1.44 0.63 1.60 1.23 ;
        RECT  1.28 1.07 2.24 1.23 ;
        RECT  2.08 1.07 2.24 1.61 ;
        RECT  2.08 1.33 2.36 1.61 ;
        RECT  1.28 1.07 1.44 2.16 ;
        RECT  0.91 2.00 1.44 2.16 ;
        RECT  0.91 2.00 1.19 2.28 ;
    END
END OR2I1SP2V1_0

MACRO OR2I1SP1V1_0
    CLASS CORE ;
    FOREIGN OR2I1SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 2.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 4.93  LAYER ME1  ;
        ANTENNADIFFAREA 2.12  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        ANTENNAMAXAREACAR 36.72  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.42 0.63 2.70 0.91 ;
        RECT  2.33 2.00 2.68 2.28 ;
        RECT  2.52 0.63 2.68 2.28 ;
        END
    END OUT
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.67 1.45 1.95 1.82 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.43 1.39 0.71 1.81 ;
        END
    END IN1
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 2.80 0.28 ;
        RECT  2.34 -0.28 2.62 0.32 ;
        RECT  1.90 0.63 2.18 0.91 ;
        RECT  1.96 -0.28 2.12 0.91 ;
        RECT  0.86 0.63 1.14 0.91 ;
        RECT  0.92 -0.28 1.08 0.91 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 2.80 3.48 ;
        RECT  2.34 2.88 2.62 3.48 ;
        RECT  1.81 2.00 2.09 2.28 ;
        RECT  1.87 2.00 2.03 3.48 ;
        RECT  0.62 2.48 0.90 2.76 ;
        RECT  0.68 2.48 0.84 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.34 0.63 0.62 0.91 ;
        RECT  0.11 0.75 0.62 0.91 ;
        RECT  0.11 1.07 1.07 1.23 ;
        RECT  0.91 1.07 1.07 1.58 ;
        RECT  0.91 1.30 1.19 1.58 ;
        RECT  0.11 0.75 0.27 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  1.35 0.63 1.66 0.91 ;
        RECT  1.35 1.07 2.36 1.23 ;
        RECT  2.08 1.07 2.36 1.35 ;
        RECT  1.35 0.63 1.51 2.16 ;
        RECT  0.91 2.00 1.51 2.16 ;
        RECT  0.91 2.00 1.19 2.28 ;
    END
END OR2I1SP1V1_0

MACRO OR2AND3SP8V1_0
    CLASS CORE ;
    FOREIGN OR2AND3SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 11.97  LAYER ME1  ;
        ANTENNADIFFAREA 6.17  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.78  LAYER ME1  ;
        ANTENNAMAXAREACAR 15.29  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.24 2.04 5.52 2.64 ;
        RECT  5.24 0.54 5.40 2.64 ;
        RECT  4.26 1.52 5.40 1.68 ;
        RECT  5.10 0.54 5.40 1.14 ;
        RECT  4.26 1.46 4.74 1.74 ;
        RECT  4.20 2.04 4.48 2.64 ;
        RECT  4.26 0.54 4.42 2.64 ;
        RECT  4.06 0.54 4.42 1.14 ;
        END
    END OUT
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.30 1.39 3.62 1.81 ;
        END
    END IN4
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.86 1.39 3.14 1.81 ;
        END
    END IN3
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 6.40 0.28 ;
        RECT  5.68 -0.28 6.22 0.32 ;
        RECT  5.62 0.54 5.90 1.14 ;
        RECT  5.68 -0.28 5.84 1.14 ;
        RECT  4.58 0.54 4.86 1.14 ;
        RECT  4.64 -0.28 4.80 1.14 ;
        RECT  3.54 0.54 3.82 1.14 ;
        RECT  3.60 -0.28 3.76 1.14 ;
        RECT  1.14 0.63 1.42 0.91 ;
        RECT  1.20 -0.28 1.36 0.91 ;
        RECT  0.10 0.63 0.38 0.91 ;
        RECT  0.16 -0.28 0.32 0.91 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 6.40 3.48 ;
        RECT  5.82 2.88 6.22 3.48 ;
        RECT  5.76 2.04 6.04 2.64 ;
        RECT  5.82 2.04 5.98 3.48 ;
        RECT  4.72 2.04 5.00 2.64 ;
        RECT  4.78 2.04 4.94 3.48 ;
        RECT  3.68 2.36 3.96 2.64 ;
        RECT  3.74 2.36 3.90 3.48 ;
        RECT  2.60 2.34 2.88 2.62 ;
        RECT  2.66 2.34 2.82 3.48 ;
        RECT  1.05 2.02 1.33 2.30 ;
        RECT  1.11 2.02 1.27 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.54 0.63 0.90 0.91 ;
        RECT  0.54 1.07 1.60 1.23 ;
        RECT  1.32 1.07 1.60 1.35 ;
        RECT  0.54 0.63 0.70 2.18 ;
        RECT  0.15 2.02 0.70 2.18 ;
        RECT  0.15 2.02 0.43 2.30 ;
        RECT  1.66 0.63 1.94 0.91 ;
        RECT  1.76 1.46 2.12 1.74 ;
        RECT  1.76 0.63 1.92 2.30 ;
        RECT  1.57 2.02 1.92 2.30 ;
        RECT  2.20 0.80 2.48 1.08 ;
        RECT  3.82 1.46 4.10 1.74 ;
        RECT  2.28 0.80 2.44 2.18 ;
        RECT  3.82 1.46 3.98 2.18 ;
        RECT  2.20 2.02 3.98 2.18 ;
        RECT  2.20 2.02 2.36 2.62 ;
        RECT  3.12 2.02 3.28 2.62 ;
        RECT  2.08 2.34 2.36 2.62 ;
        RECT  3.12 2.34 3.40 2.62 ;
    END
END OR2AND3SP8V1_0

MACRO OR2AND3SP4V1_0
    CLASS CORE ;
    FOREIGN OR2AND3SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.86 1.39 3.14 1.81 ;
        END
    END IN3
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.30 1.39 3.62 1.81 ;
        END
    END IN4
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 9.61  LAYER ME1  ;
        ANTENNADIFFAREA 4.62  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER ME1  ;
        ANTENNAMAXAREACAR 19.44  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.26 1.46 4.72 1.74 ;
        RECT  4.20 2.04 4.48 2.64 ;
        RECT  4.26 0.54 4.42 2.64 ;
        RECT  4.06 0.54 4.42 1.14 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 5.20 3.48 ;
        RECT  4.74 2.88 5.02 3.48 ;
        RECT  4.72 2.04 5.00 2.64 ;
        RECT  4.78 2.04 4.94 3.48 ;
        RECT  3.68 2.36 3.96 2.64 ;
        RECT  3.74 2.36 3.90 3.48 ;
        RECT  2.60 2.34 2.88 2.62 ;
        RECT  2.66 2.34 2.82 3.48 ;
        RECT  1.05 2.02 1.33 2.30 ;
        RECT  1.11 2.02 1.27 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 5.20 0.28 ;
        RECT  4.64 -0.28 5.02 0.32 ;
        RECT  4.58 0.54 4.86 1.14 ;
        RECT  4.64 -0.28 4.80 1.14 ;
        RECT  3.54 0.54 3.82 1.14 ;
        RECT  3.60 -0.28 3.76 1.14 ;
        RECT  1.14 0.63 1.42 0.91 ;
        RECT  1.20 -0.28 1.36 0.91 ;
        RECT  0.10 0.63 0.38 0.91 ;
        RECT  0.16 -0.28 0.32 0.91 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.54 0.63 0.90 0.91 ;
        RECT  0.54 1.07 1.60 1.23 ;
        RECT  1.32 1.07 1.60 1.35 ;
        RECT  0.54 0.63 0.70 2.18 ;
        RECT  0.15 2.02 0.70 2.18 ;
        RECT  0.15 2.02 0.43 2.30 ;
        RECT  1.66 0.63 1.94 0.91 ;
        RECT  1.76 1.46 2.12 1.74 ;
        RECT  1.76 0.63 1.92 2.30 ;
        RECT  1.57 2.02 1.92 2.30 ;
        RECT  2.20 0.80 2.48 1.08 ;
        RECT  3.82 1.46 4.10 1.74 ;
        RECT  2.28 0.80 2.44 2.18 ;
        RECT  3.82 1.46 3.98 2.18 ;
        RECT  2.20 2.02 3.98 2.18 ;
        RECT  2.20 2.02 2.36 2.62 ;
        RECT  3.12 2.02 3.28 2.62 ;
        RECT  2.08 2.34 2.36 2.62 ;
        RECT  3.12 2.34 3.40 2.62 ;
    END
END OR2AND3SP4V1_0

MACRO OR2AND3SP2V1_0
    CLASS CORE ;
    FOREIGN OR2AND3SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 8.67  LAYER ME1  ;
        ANTENNADIFFAREA 4.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.28  LAYER ME1  ;
        ANTENNAMAXAREACAR 31.15  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.26 1.46 4.72 1.74 ;
        RECT  4.20 2.06 4.48 2.34 ;
        RECT  4.26 0.54 4.42 2.34 ;
        RECT  4.04 0.54 4.42 1.14 ;
        END
    END OUT
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.30 1.39 3.62 1.81 ;
        END
    END IN4
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.86 1.39 3.14 1.81 ;
        END
    END IN3
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.80 0.28 ;
        RECT  4.34 -0.28 4.62 0.32 ;
        RECT  3.52 0.54 3.80 1.14 ;
        RECT  3.58 -0.28 3.74 1.14 ;
        RECT  1.14 0.63 1.42 0.91 ;
        RECT  1.20 -0.28 1.36 0.91 ;
        RECT  0.10 0.63 0.38 0.91 ;
        RECT  0.16 -0.28 0.32 0.91 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.80 3.48 ;
        RECT  4.34 2.88 4.62 3.48 ;
        RECT  3.68 2.38 3.96 2.66 ;
        RECT  3.74 2.38 3.90 3.48 ;
        RECT  2.60 2.34 2.88 2.62 ;
        RECT  2.66 2.34 2.82 3.48 ;
        RECT  1.05 2.02 1.33 2.30 ;
        RECT  1.11 2.02 1.27 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.54 0.63 0.90 0.91 ;
        RECT  0.54 1.07 1.60 1.23 ;
        RECT  1.32 1.07 1.60 1.35 ;
        RECT  0.54 0.63 0.70 2.18 ;
        RECT  0.15 2.02 0.70 2.18 ;
        RECT  0.15 2.02 0.43 2.30 ;
        RECT  1.66 0.63 1.94 0.91 ;
        RECT  1.76 1.46 2.12 1.74 ;
        RECT  1.76 0.63 1.92 2.30 ;
        RECT  1.57 2.02 1.92 2.30 ;
        RECT  2.20 0.80 2.48 1.08 ;
        RECT  3.82 1.46 4.10 1.74 ;
        RECT  2.28 0.80 2.44 2.18 ;
        RECT  3.82 1.46 3.98 2.18 ;
        RECT  2.20 2.02 3.98 2.18 ;
        RECT  2.20 2.02 2.36 2.62 ;
        RECT  3.12 2.02 3.28 2.62 ;
        RECT  2.08 2.34 2.36 2.62 ;
        RECT  3.12 2.34 3.40 2.62 ;
    END
END OR2AND3SP2V1_0

MACRO OR2AND3SP1V1_0
    CLASS CORE ;
    FOREIGN OR2AND3SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.30 1.39 3.62 1.81 ;
        END
    END IN4
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 8.50  LAYER ME1  ;
        ANTENNADIFFAREA 3.55  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        ANTENNAMAXAREACAR 42.18  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.26 1.46 4.72 1.74 ;
        RECT  4.16 2.34 4.44 2.62 ;
        RECT  4.26 0.80 4.42 2.62 ;
        RECT  4.00 0.80 4.42 1.08 ;
        END
    END OUT
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.86 1.39 3.14 1.81 ;
        END
    END IN3
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.80 0.28 ;
        RECT  4.34 -0.28 4.62 0.32 ;
        RECT  3.48 0.80 3.76 1.08 ;
        RECT  3.52 -0.28 3.68 1.08 ;
        RECT  1.14 0.63 1.42 0.91 ;
        RECT  1.20 -0.28 1.36 0.91 ;
        RECT  0.10 0.63 0.38 0.91 ;
        RECT  0.16 -0.28 0.32 0.91 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.80 3.48 ;
        RECT  4.34 2.88 4.62 3.48 ;
        RECT  3.64 2.34 3.92 2.62 ;
        RECT  3.70 2.34 3.86 3.48 ;
        RECT  2.60 2.34 2.88 2.62 ;
        RECT  2.66 2.34 2.82 3.48 ;
        RECT  1.05 2.02 1.33 2.30 ;
        RECT  1.11 2.02 1.27 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.54 0.63 0.90 0.91 ;
        RECT  0.54 1.07 1.60 1.23 ;
        RECT  1.32 1.07 1.60 1.35 ;
        RECT  0.54 0.63 0.70 2.18 ;
        RECT  0.15 2.02 0.70 2.18 ;
        RECT  0.15 2.02 0.43 2.30 ;
        RECT  1.66 0.63 1.94 0.91 ;
        RECT  1.76 1.46 2.12 1.74 ;
        RECT  1.76 0.63 1.92 2.30 ;
        RECT  1.57 2.02 1.92 2.30 ;
        RECT  2.20 0.80 2.48 1.08 ;
        RECT  2.28 0.80 2.44 2.18 ;
        RECT  3.82 1.90 4.10 2.18 ;
        RECT  2.20 2.02 4.10 2.18 ;
        RECT  2.20 2.02 2.36 2.62 ;
        RECT  3.12 2.02 3.28 2.62 ;
        RECT  2.08 2.34 2.36 2.62 ;
        RECT  3.12 2.34 3.40 2.62 ;
    END
END OR2AND3SP1V1_0

MACRO OR2AND2SP8V1_0
    CLASS CORE ;
    FOREIGN OR2AND2SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 10.87  LAYER ME1  ;
        ANTENNADIFFAREA 5.99  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.71  LAYER ME1  ;
        ANTENNAMAXAREACAR 15.31  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.70 1.97 4.98 2.57 ;
        RECT  4.70 0.63 4.98 1.23 ;
        RECT  4.70 0.63 4.86 2.57 ;
        RECT  3.78 1.52 4.86 1.68 ;
        RECT  3.66 1.97 3.94 2.57 ;
        RECT  3.78 0.63 3.94 2.57 ;
        RECT  3.66 0.63 3.94 1.23 ;
        END
    END OUT
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.86 1.39 3.14 1.81 ;
        END
    END IN3
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 5.60 3.48 ;
        RECT  5.22 1.97 5.50 2.57 ;
        RECT  5.14 2.88 5.44 3.48 ;
        RECT  5.28 1.97 5.44 3.48 ;
        RECT  4.18 1.97 4.46 2.57 ;
        RECT  4.24 1.97 4.40 3.48 ;
        RECT  3.14 1.97 3.42 2.57 ;
        RECT  3.20 1.97 3.36 3.48 ;
        RECT  2.02 1.97 2.30 2.25 ;
        RECT  2.12 1.97 2.28 3.48 ;
        RECT  1.00 2.02 1.28 2.30 ;
        RECT  1.11 2.02 1.27 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 5.60 0.28 ;
        RECT  5.22 0.63 5.50 1.23 ;
        RECT  5.28 -0.28 5.44 1.23 ;
        RECT  5.14 -0.28 5.44 0.32 ;
        RECT  4.18 0.63 4.46 1.23 ;
        RECT  4.24 -0.28 4.40 1.23 ;
        RECT  3.14 0.63 3.42 0.91 ;
        RECT  3.20 -0.28 3.36 0.91 ;
        RECT  1.14 0.63 1.42 0.91 ;
        RECT  1.20 -0.28 1.36 0.91 ;
        RECT  0.10 0.63 0.38 0.91 ;
        RECT  0.16 -0.28 0.32 0.91 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.54 0.63 0.90 0.91 ;
        RECT  0.54 1.07 1.58 1.23 ;
        RECT  1.30 1.07 1.58 1.35 ;
        RECT  0.54 0.63 0.70 2.18 ;
        RECT  0.10 2.02 0.70 2.18 ;
        RECT  0.10 2.02 0.38 2.30 ;
        RECT  1.66 0.63 1.94 0.91 ;
        RECT  1.74 0.63 1.90 1.68 ;
        RECT  1.64 1.52 2.34 1.68 ;
        RECT  2.06 1.46 2.34 1.74 ;
        RECT  1.64 1.52 1.80 2.30 ;
        RECT  1.52 2.02 1.80 2.30 ;
        RECT  2.20 0.63 2.66 0.91 ;
        RECT  2.50 1.07 3.50 1.23 ;
        RECT  3.34 1.07 3.50 1.67 ;
        RECT  3.34 1.39 3.62 1.67 ;
        RECT  2.50 0.63 2.66 2.25 ;
        RECT  2.50 1.97 2.86 2.25 ;
    END
END OR2AND2SP8V1_0

MACRO OR2AND2SP4V1_0
    CLASS CORE ;
    FOREIGN OR2AND2SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 9.04  LAYER ME1  ;
        ANTENNADIFFAREA 4.54  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.42  LAYER ME1  ;
        ANTENNAMAXAREACAR 21.39  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.78 1.52 4.28 1.68 ;
        RECT  3.70 1.97 3.98 2.57 ;
        RECT  3.78 0.63 3.94 2.57 ;
        RECT  3.66 0.63 3.94 1.23 ;
        END
    END OUT
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.86 1.39 3.14 1.81 ;
        END
    END IN3
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.80 0.28 ;
        RECT  4.24 -0.28 4.62 0.32 ;
        RECT  4.18 0.63 4.46 1.23 ;
        RECT  4.24 -0.28 4.40 1.23 ;
        RECT  3.14 0.63 3.42 0.91 ;
        RECT  3.20 -0.28 3.36 0.91 ;
        RECT  1.14 0.63 1.42 0.91 ;
        RECT  1.20 -0.28 1.36 0.91 ;
        RECT  0.10 0.63 0.38 0.91 ;
        RECT  0.16 -0.28 0.32 0.91 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.80 3.48 ;
        RECT  4.28 2.88 4.62 3.48 ;
        RECT  4.22 1.97 4.50 2.57 ;
        RECT  4.28 1.97 4.44 3.48 ;
        RECT  3.18 1.97 3.46 2.57 ;
        RECT  3.24 1.97 3.40 3.48 ;
        RECT  2.06 1.97 2.34 2.25 ;
        RECT  2.12 1.97 2.28 3.48 ;
        RECT  1.00 2.02 1.28 2.30 ;
        RECT  1.11 2.02 1.27 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.54 0.63 0.90 0.91 ;
        RECT  0.54 1.07 1.58 1.23 ;
        RECT  1.30 1.07 1.58 1.35 ;
        RECT  0.54 0.63 0.70 2.18 ;
        RECT  0.10 2.02 0.70 2.18 ;
        RECT  0.10 2.02 0.38 2.30 ;
        RECT  1.66 0.63 1.94 0.91 ;
        RECT  1.74 1.52 2.34 1.68 ;
        RECT  2.06 1.46 2.34 1.74 ;
        RECT  1.74 0.63 1.90 2.30 ;
        RECT  1.52 2.02 1.90 2.30 ;
        RECT  2.20 0.63 2.66 0.91 ;
        RECT  2.50 1.07 3.50 1.23 ;
        RECT  3.34 1.07 3.50 1.67 ;
        RECT  3.34 1.39 3.62 1.67 ;
        RECT  2.50 0.63 2.66 2.25 ;
        RECT  2.50 1.97 2.90 2.25 ;
    END
END OR2AND2SP4V1_0

MACRO OR2AND2SP2V1_0
    CLASS CORE ;
    FOREIGN OR2AND2SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 7.18  LAYER ME1  ;
        ANTENNADIFFAREA 3.59  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.28  LAYER ME1  ;
        ANTENNAMAXAREACAR 25.78  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.62 2.00 3.90 2.60 ;
        RECT  3.62 0.63 3.90 1.23 ;
        RECT  3.72 0.63 3.88 2.60 ;
        END
    END OUT
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.80 1.39 3.12 1.81 ;
        END
    END IN3
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.00 0.28 ;
        RECT  3.54 -0.28 3.82 0.32 ;
        RECT  3.10 0.63 3.38 0.91 ;
        RECT  3.16 -0.28 3.32 0.91 ;
        RECT  1.14 0.63 1.42 0.91 ;
        RECT  1.20 -0.28 1.36 0.91 ;
        RECT  0.10 0.63 0.38 0.91 ;
        RECT  0.16 -0.28 0.32 0.91 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.00 3.48 ;
        RECT  3.54 2.88 3.82 3.48 ;
        RECT  3.10 2.00 3.38 2.60 ;
        RECT  3.16 2.00 3.32 3.48 ;
        RECT  1.98 2.47 2.26 2.75 ;
        RECT  2.04 2.47 2.20 3.48 ;
        RECT  1.00 2.00 1.28 2.28 ;
        RECT  1.07 2.00 1.23 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.54 0.63 0.90 0.91 ;
        RECT  0.54 1.07 1.58 1.23 ;
        RECT  1.30 1.07 1.58 1.35 ;
        RECT  0.54 0.63 0.70 2.16 ;
        RECT  0.10 2.00 0.70 2.16 ;
        RECT  0.10 2.00 0.38 2.28 ;
        RECT  1.66 0.63 1.94 0.91 ;
        RECT  1.78 1.54 2.32 1.82 ;
        RECT  1.78 0.63 1.94 2.28 ;
        RECT  1.52 2.00 1.94 2.28 ;
        RECT  2.16 0.63 2.64 0.91 ;
        RECT  2.48 1.07 3.44 1.23 ;
        RECT  3.28 1.07 3.44 1.66 ;
        RECT  3.28 1.38 3.56 1.66 ;
        RECT  2.48 0.63 2.64 2.75 ;
        RECT  2.48 2.47 2.82 2.75 ;
    END
END OR2AND2SP2V1_0

MACRO OR2AND2SP1V1_0
    CLASS CORE ;
    FOREIGN OR2AND2SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 7.08  LAYER ME1  ;
        ANTENNADIFFAREA 3.09  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        ANTENNAMAXAREACAR 35.14  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.62 1.97 3.91 2.25 ;
        RECT  3.75 0.63 3.91 2.25 ;
        RECT  3.72 1.52 3.91 1.68 ;
        RECT  3.62 0.63 3.91 0.91 ;
        END
    END OUT
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.86 1.39 3.14 1.81 ;
        END
    END IN3
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.00 0.28 ;
        RECT  3.54 -0.28 3.82 0.32 ;
        RECT  3.10 0.63 3.38 0.91 ;
        RECT  3.16 -0.28 3.32 0.91 ;
        RECT  1.14 0.63 1.42 0.91 ;
        RECT  1.20 -0.28 1.36 0.91 ;
        RECT  0.10 0.63 0.38 0.91 ;
        RECT  0.16 -0.28 0.32 0.91 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.00 3.48 ;
        RECT  3.54 2.88 3.82 3.48 ;
        RECT  3.10 1.97 3.38 2.25 ;
        RECT  3.16 1.97 3.32 3.48 ;
        RECT  2.06 1.97 2.34 2.25 ;
        RECT  2.12 1.97 2.28 3.48 ;
        RECT  1.00 2.02 1.28 2.30 ;
        RECT  1.11 2.02 1.27 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.54 0.63 0.90 0.91 ;
        RECT  0.54 1.07 1.58 1.23 ;
        RECT  1.30 1.07 1.58 1.35 ;
        RECT  0.54 0.63 0.70 2.18 ;
        RECT  0.10 2.02 0.70 2.18 ;
        RECT  0.10 2.02 0.38 2.30 ;
        RECT  1.66 0.63 1.94 0.91 ;
        RECT  1.74 1.52 2.34 1.68 ;
        RECT  2.06 1.46 2.34 1.74 ;
        RECT  1.74 0.63 1.90 2.30 ;
        RECT  1.52 2.02 1.90 2.30 ;
        RECT  2.20 0.63 2.66 0.91 ;
        RECT  2.50 1.07 3.59 1.23 ;
        RECT  3.31 1.07 3.59 1.35 ;
        RECT  2.50 0.63 2.66 2.25 ;
        RECT  2.50 1.97 2.86 2.25 ;
    END
END OR2AND2SP1V1_0

MACRO OR23NAND3SP8V1_0
    CLASS CORE ;
    FOREIGN OR23NAND3SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 14.94  LAYER ME1  ;
        ANTENNADIFFAREA 7.59  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.78  LAYER ME1  ;
        ANTENNAMAXAREACAR 19.21  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.84 0.63 7.14 1.23 ;
        RECT  6.72 1.92 7.00 2.52 ;
        RECT  6.84 0.63 7.00 2.52 ;
        RECT  5.84 1.52 7.00 1.68 ;
        RECT  5.84 1.46 6.32 1.74 ;
        RECT  5.82 0.63 6.10 1.23 ;
        RECT  5.68 1.92 6.00 2.52 ;
        RECT  5.84 0.63 6.00 2.52 ;
        END
    END OUT
    PIN IN6
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.26 0.99 3.54 1.41 ;
        END
    END IN6
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.36 1.62 1.81 ;
        END
    END IN3
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.10 1.47 2.51 1.76 ;
        RECT  2.10 1.47 2.38 1.78 ;
        END
    END IN4
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN5
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.41 0.97 2.74 1.31 ;
        END
    END IN5
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 8.00 3.48 ;
        RECT  7.30 2.88 7.82 3.48 ;
        RECT  7.24 1.92 7.52 2.52 ;
        RECT  7.30 1.92 7.46 3.48 ;
        RECT  6.20 1.92 6.48 2.52 ;
        RECT  6.26 1.92 6.42 3.48 ;
        RECT  5.16 1.92 5.44 2.52 ;
        RECT  5.22 1.92 5.38 3.48 ;
        RECT  3.36 1.92 3.64 2.20 ;
        RECT  3.42 1.92 3.58 3.48 ;
        RECT  1.08 2.02 1.36 2.30 ;
        RECT  1.14 2.02 1.30 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 8.00 0.28 ;
        RECT  7.44 -0.28 7.82 0.32 ;
        RECT  7.38 0.63 7.66 1.23 ;
        RECT  7.44 -0.28 7.60 1.23 ;
        RECT  6.34 0.63 6.62 1.23 ;
        RECT  6.40 -0.28 6.56 1.23 ;
        RECT  5.30 0.63 5.58 1.23 ;
        RECT  5.36 -0.28 5.52 1.23 ;
        RECT  4.22 0.63 4.50 0.91 ;
        RECT  4.28 -0.28 4.44 0.91 ;
        RECT  3.22 0.53 3.50 0.81 ;
        RECT  3.28 -0.28 3.44 0.81 ;
        RECT  2.18 0.53 2.46 0.81 ;
        RECT  2.24 -0.28 2.40 0.81 ;
        RECT  1.14 0.53 1.42 0.81 ;
        RECT  1.20 -0.28 1.36 0.81 ;
        RECT  0.10 0.53 0.38 0.81 ;
        RECT  0.16 -0.28 0.32 0.81 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.54 0.53 0.90 0.81 ;
        RECT  0.54 0.53 0.70 2.18 ;
        RECT  0.22 2.02 0.70 2.18 ;
        RECT  0.22 2.02 0.52 2.30 ;
        RECT  0.22 2.02 0.38 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  1.66 0.53 1.94 0.81 ;
        RECT  1.78 0.53 1.94 2.30 ;
        RECT  1.78 2.02 2.20 2.30 ;
        RECT  2.04 2.02 2.20 2.70 ;
        RECT  2.04 2.42 2.34 2.70 ;
        RECT  2.70 0.53 3.06 0.81 ;
        RECT  4.02 1.48 4.30 1.76 ;
        RECT  2.90 1.60 4.30 1.76 ;
        RECT  2.90 0.53 3.06 2.08 ;
        RECT  2.46 1.92 3.06 2.08 ;
        RECT  2.46 1.92 2.74 2.20 ;
        RECT  3.70 0.63 3.98 0.91 ;
        RECT  4.74 0.63 5.02 0.91 ;
        RECT  3.82 0.63 3.98 1.32 ;
        RECT  3.82 1.16 4.62 1.32 ;
        RECT  4.80 0.63 4.96 1.55 ;
        RECT  4.46 1.39 5.68 1.55 ;
        RECT  5.40 1.39 5.68 1.67 ;
        RECT  4.46 1.16 4.62 2.08 ;
        RECT  3.84 1.92 4.62 2.08 ;
        RECT  3.84 1.92 4.12 2.20 ;
    END
END OR23NAND3SP8V1_0

MACRO OR23NAND3SP4V1_0
    CLASS CORE ;
    FOREIGN OR23NAND3SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN5
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.41 0.97 2.74 1.31 ;
        END
    END IN5
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.10 1.47 2.51 1.76 ;
        RECT  2.10 1.47 2.38 1.78 ;
        END
    END IN4
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.36 1.62 1.81 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN IN6
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.26 0.99 3.54 1.41 ;
        END
    END IN6
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 12.59  LAYER ME1  ;
        ANTENNADIFFAREA 5.88  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER ME1  ;
        ANTENNAMAXAREACAR 25.71  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.84 1.46 6.32 1.74 ;
        RECT  5.82 0.63 6.10 1.23 ;
        RECT  5.68 1.92 6.00 2.52 ;
        RECT  5.84 0.63 6.00 2.52 ;
        END
    END OUT
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 6.80 0.28 ;
        RECT  6.34 0.63 6.62 1.23 ;
        RECT  6.34 -0.28 6.62 0.32 ;
        RECT  6.40 -0.28 6.56 1.23 ;
        RECT  5.30 0.63 5.58 1.23 ;
        RECT  5.36 -0.28 5.52 1.23 ;
        RECT  4.22 0.63 4.50 0.91 ;
        RECT  4.28 -0.28 4.44 0.91 ;
        RECT  3.22 0.53 3.50 0.81 ;
        RECT  3.28 -0.28 3.44 0.81 ;
        RECT  2.18 0.53 2.46 0.81 ;
        RECT  2.24 -0.28 2.40 0.81 ;
        RECT  1.14 0.53 1.42 0.81 ;
        RECT  1.20 -0.28 1.36 0.81 ;
        RECT  0.10 0.53 0.38 0.81 ;
        RECT  0.16 -0.28 0.32 0.81 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 6.80 3.48 ;
        RECT  6.26 2.88 6.62 3.48 ;
        RECT  6.20 1.92 6.48 2.52 ;
        RECT  6.26 1.92 6.42 3.48 ;
        RECT  5.16 1.92 5.44 2.52 ;
        RECT  5.22 1.92 5.38 3.48 ;
        RECT  3.36 1.92 3.64 2.20 ;
        RECT  3.42 1.92 3.58 3.48 ;
        RECT  1.08 2.02 1.36 2.30 ;
        RECT  1.14 2.02 1.30 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.54 0.53 0.90 0.81 ;
        RECT  0.54 0.53 0.70 2.18 ;
        RECT  0.22 2.02 0.70 2.18 ;
        RECT  0.22 2.02 0.52 2.30 ;
        RECT  0.22 2.02 0.38 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  1.66 0.53 1.94 0.81 ;
        RECT  1.78 0.53 1.94 2.30 ;
        RECT  1.78 2.02 2.20 2.30 ;
        RECT  2.04 2.02 2.20 2.70 ;
        RECT  2.04 2.42 2.34 2.70 ;
        RECT  2.70 0.53 3.06 0.81 ;
        RECT  4.02 1.48 4.30 1.76 ;
        RECT  2.90 1.60 4.30 1.76 ;
        RECT  2.90 0.53 3.06 2.08 ;
        RECT  2.46 1.92 3.06 2.08 ;
        RECT  2.46 1.92 2.74 2.20 ;
        RECT  3.70 0.63 3.98 0.91 ;
        RECT  4.74 0.63 5.02 0.91 ;
        RECT  3.82 0.63 3.98 1.32 ;
        RECT  3.82 1.16 4.62 1.32 ;
        RECT  4.80 0.63 4.96 1.55 ;
        RECT  4.46 1.39 5.68 1.55 ;
        RECT  5.40 1.39 5.68 1.67 ;
        RECT  4.46 1.16 4.62 2.08 ;
        RECT  3.84 1.92 4.62 2.08 ;
        RECT  3.84 1.92 4.12 2.20 ;
    END
END OR23NAND3SP4V1_0

MACRO OR23NAND3SP2V1_0
    CLASS CORE ;
    FOREIGN OR23NAND3SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 11.69  LAYER ME1  ;
        ANTENNADIFFAREA 5.15  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.35  LAYER ME1  ;
        ANTENNAMAXAREACAR 33.83  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.84 1.46 6.32 1.74 ;
        RECT  5.82 0.63 6.10 1.23 ;
        RECT  5.68 1.92 6.00 2.52 ;
        RECT  5.84 0.63 6.00 2.52 ;
        END
    END OUT
    PIN IN6
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.26 0.99 3.54 1.41 ;
        END
    END IN6
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.36 1.62 1.81 ;
        END
    END IN3
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.10 1.47 2.51 1.76 ;
        RECT  2.10 1.47 2.38 1.78 ;
        END
    END IN4
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN5
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.41 0.97 2.74 1.31 ;
        END
    END IN5
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 6.40 3.48 ;
        RECT  5.94 2.88 6.22 3.48 ;
        RECT  5.16 1.92 5.44 2.52 ;
        RECT  5.22 1.92 5.38 3.48 ;
        RECT  3.36 1.92 3.64 2.20 ;
        RECT  3.42 1.92 3.58 3.48 ;
        RECT  1.08 2.02 1.36 2.30 ;
        RECT  1.14 2.02 1.30 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 6.40 0.28 ;
        RECT  5.94 -0.28 6.22 0.32 ;
        RECT  5.30 0.63 5.58 1.23 ;
        RECT  5.36 -0.28 5.52 1.23 ;
        RECT  4.22 0.63 4.50 0.91 ;
        RECT  4.28 -0.28 4.44 0.91 ;
        RECT  3.22 0.53 3.50 0.81 ;
        RECT  3.28 -0.28 3.44 0.81 ;
        RECT  2.18 0.53 2.46 0.81 ;
        RECT  2.24 -0.28 2.40 0.81 ;
        RECT  1.14 0.53 1.42 0.81 ;
        RECT  1.20 -0.28 1.36 0.81 ;
        RECT  0.10 0.53 0.38 0.81 ;
        RECT  0.16 -0.28 0.32 0.81 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.54 0.53 0.90 0.81 ;
        RECT  0.54 0.53 0.70 2.18 ;
        RECT  0.22 2.02 0.70 2.18 ;
        RECT  0.22 2.02 0.52 2.30 ;
        RECT  0.22 2.02 0.38 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  1.66 0.53 1.94 0.81 ;
        RECT  1.78 0.53 1.94 2.30 ;
        RECT  1.78 2.02 2.20 2.30 ;
        RECT  2.04 2.02 2.20 2.70 ;
        RECT  2.04 2.42 2.34 2.70 ;
        RECT  2.70 0.53 3.06 0.81 ;
        RECT  4.02 1.48 4.30 1.76 ;
        RECT  2.90 1.60 4.30 1.76 ;
        RECT  2.90 0.53 3.06 2.08 ;
        RECT  2.46 1.92 3.06 2.08 ;
        RECT  2.46 1.92 2.74 2.20 ;
        RECT  3.70 0.63 3.98 0.91 ;
        RECT  4.74 0.63 5.02 0.91 ;
        RECT  3.82 0.63 3.98 1.32 ;
        RECT  3.82 1.16 4.62 1.32 ;
        RECT  4.80 0.63 4.96 1.55 ;
        RECT  4.46 1.39 5.68 1.55 ;
        RECT  5.40 1.39 5.68 1.67 ;
        RECT  4.46 1.16 4.62 2.08 ;
        RECT  3.84 1.92 4.62 2.08 ;
        RECT  3.84 1.92 4.12 2.20 ;
    END
END OR23NAND3SP2V1_0

MACRO OR23NAND3SP1V1_0
    CLASS CORE ;
    FOREIGN OR23NAND3SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 10.97  LAYER ME1  ;
        ANTENNADIFFAREA 4.70  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.27  LAYER ME1  ;
        ANTENNAMAXAREACAR 40.80  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.84 1.46 6.32 1.74 ;
        RECT  5.78 0.63 6.06 0.91 ;
        RECT  5.64 1.92 6.00 2.20 ;
        RECT  5.84 0.63 6.00 2.20 ;
        END
    END OUT
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.36 1.62 1.81 ;
        END
    END IN3
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.10 1.47 2.51 1.76 ;
        RECT  2.10 1.47 2.38 1.78 ;
        END
    END IN4
    PIN IN5
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.41 0.97 2.74 1.31 ;
        END
    END IN5
    PIN IN6
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.26 0.99 3.54 1.41 ;
        END
    END IN6
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 6.40 3.48 ;
        RECT  5.94 2.88 6.22 3.48 ;
        RECT  5.12 1.92 5.40 2.20 ;
        RECT  5.18 1.92 5.34 3.48 ;
        RECT  3.36 1.92 3.64 2.20 ;
        RECT  3.42 1.92 3.58 3.48 ;
        RECT  1.08 2.02 1.36 2.30 ;
        RECT  1.14 2.02 1.30 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 6.40 0.28 ;
        RECT  5.94 -0.28 6.22 0.32 ;
        RECT  5.26 0.63 5.54 0.91 ;
        RECT  5.32 -0.28 5.48 0.91 ;
        RECT  4.22 0.63 4.50 0.91 ;
        RECT  4.28 -0.28 4.44 0.91 ;
        RECT  3.22 0.53 3.50 0.81 ;
        RECT  3.28 -0.28 3.44 0.81 ;
        RECT  2.18 0.53 2.46 0.81 ;
        RECT  2.24 -0.28 2.40 0.81 ;
        RECT  1.14 0.53 1.42 0.81 ;
        RECT  1.20 -0.28 1.36 0.81 ;
        RECT  0.10 0.53 0.38 0.81 ;
        RECT  0.16 -0.28 0.32 0.81 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.54 0.53 0.90 0.81 ;
        RECT  0.54 0.53 0.70 2.18 ;
        RECT  0.22 2.02 0.70 2.18 ;
        RECT  0.22 2.02 0.52 2.30 ;
        RECT  0.22 2.02 0.38 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  1.66 0.53 1.94 0.81 ;
        RECT  1.78 0.53 1.94 2.30 ;
        RECT  1.78 2.02 2.20 2.30 ;
        RECT  2.04 2.02 2.20 2.70 ;
        RECT  2.04 2.42 2.34 2.70 ;
        RECT  2.70 0.53 3.06 0.81 ;
        RECT  4.02 1.48 4.30 1.76 ;
        RECT  2.90 1.60 4.30 1.76 ;
        RECT  2.90 0.53 3.06 2.08 ;
        RECT  2.46 1.92 3.06 2.08 ;
        RECT  2.46 1.92 2.74 2.20 ;
        RECT  3.70 0.63 3.98 0.91 ;
        RECT  4.74 0.63 5.02 0.91 ;
        RECT  3.82 0.63 3.98 1.32 ;
        RECT  4.80 0.63 4.96 1.32 ;
        RECT  3.82 1.16 5.68 1.32 ;
        RECT  5.40 1.10 5.68 1.38 ;
        RECT  4.46 1.16 4.62 2.08 ;
        RECT  3.84 1.92 4.62 2.08 ;
        RECT  3.84 1.92 4.12 2.20 ;
    END
END OR23NAND3SP1V1_0

MACRO OR23AND3SP8V1_0
    CLASS CORE ;
    FOREIGN OR23AND3SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 16.30  LAYER ME1  ;
        ANTENNADIFFAREA 8.85  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.95  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.23  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.58 1.84 7.86 2.44 ;
        RECT  7.58 0.64 7.86 1.24 ;
        RECT  7.58 0.64 7.74 2.44 ;
        RECT  6.66 1.52 7.74 1.68 ;
        RECT  6.54 1.84 6.82 2.44 ;
        RECT  6.66 0.64 6.82 2.44 ;
        RECT  6.54 0.64 6.82 1.24 ;
        END
    END OUT
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.39 1.62 1.81 ;
        END
    END IN3
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.10 1.39 2.38 1.81 ;
        END
    END IN4
    PIN IN5
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.86 1.39 3.14 1.76 ;
        END
    END IN5
    PIN IN6
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.30 1.39 3.62 1.76 ;
        END
    END IN6
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 8.80 0.28 ;
        RECT  8.34 -0.28 8.62 0.32 ;
        RECT  8.10 0.64 8.38 1.24 ;
        RECT  8.16 -0.28 8.32 1.24 ;
        RECT  7.06 0.64 7.34 1.24 ;
        RECT  7.12 -0.28 7.28 1.24 ;
        RECT  5.98 0.54 6.26 1.24 ;
        RECT  6.04 -0.28 6.20 1.24 ;
        RECT  4.46 0.63 4.74 0.91 ;
        RECT  4.52 -0.28 4.68 0.91 ;
        RECT  3.42 0.63 3.70 0.91 ;
        RECT  3.48 -0.28 3.64 0.91 ;
        RECT  2.28 0.63 2.56 0.91 ;
        RECT  2.34 -0.28 2.50 0.91 ;
        RECT  1.14 0.63 1.42 0.91 ;
        RECT  1.20 -0.28 1.36 0.91 ;
        RECT  0.10 0.63 0.38 0.91 ;
        RECT  0.16 -0.28 0.32 0.91 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 8.80 3.48 ;
        RECT  8.18 2.88 8.62 3.48 ;
        RECT  8.10 1.84 8.38 2.44 ;
        RECT  8.18 1.84 8.34 3.48 ;
        RECT  7.06 1.84 7.34 2.44 ;
        RECT  7.12 1.84 7.28 3.48 ;
        RECT  5.98 1.84 6.26 2.54 ;
        RECT  6.04 1.84 6.20 3.48 ;
        RECT  3.58 1.92 3.86 2.20 ;
        RECT  3.64 1.92 3.80 3.48 ;
        RECT  1.14 2.02 1.42 2.30 ;
        RECT  1.20 2.02 1.36 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.54 0.63 0.90 0.91 ;
        RECT  0.54 0.63 0.70 2.18 ;
        RECT  0.24 2.02 0.70 2.18 ;
        RECT  0.24 2.02 0.52 2.30 ;
        RECT  0.24 2.02 0.40 2.76 ;
        RECT  0.10 2.48 0.40 2.76 ;
        RECT  1.66 0.63 1.94 0.91 ;
        RECT  1.78 0.63 1.94 2.18 ;
        RECT  1.78 2.02 2.32 2.18 ;
        RECT  2.04 2.02 2.32 2.30 ;
        RECT  2.16 2.02 2.32 2.70 ;
        RECT  2.16 2.42 2.46 2.70 ;
        RECT  2.90 0.63 3.18 0.91 ;
        RECT  2.90 0.63 3.06 1.23 ;
        RECT  2.54 1.07 3.98 1.23 ;
        RECT  3.82 1.07 3.98 1.74 ;
        RECT  3.82 1.46 4.10 1.74 ;
        RECT  2.54 1.07 2.70 2.20 ;
        RECT  2.54 1.92 2.96 2.20 ;
        RECT  3.94 0.63 4.30 0.91 ;
        RECT  4.98 0.63 5.26 0.91 ;
        RECT  4.14 0.63 4.30 1.23 ;
        RECT  4.14 1.07 5.14 1.23 ;
        RECT  4.98 1.40 5.42 1.68 ;
        RECT  4.98 0.63 5.14 2.20 ;
        RECT  4.86 1.92 5.14 2.20 ;
        RECT  5.46 0.54 5.74 1.24 ;
        RECT  5.58 1.46 6.48 1.62 ;
        RECT  6.20 1.40 6.48 1.68 ;
        RECT  5.58 0.54 5.74 2.54 ;
        RECT  5.46 1.84 5.74 2.54 ;
    END
END OR23AND3SP8V1_0

MACRO OR23AND3SP4V1_0
    CLASS CORE ;
    FOREIGN OR23AND3SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 13.37  LAYER ME1  ;
        ANTENNADIFFAREA 6.82  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.62  LAYER ME1  ;
        ANTENNAMAXAREACAR 21.59  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.66 1.52 7.08 1.68 ;
        RECT  6.54 1.84 6.82 2.44 ;
        RECT  6.66 0.64 6.82 2.44 ;
        RECT  6.54 0.64 6.82 1.24 ;
        END
    END OUT
    PIN IN6
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.30 1.39 3.62 1.76 ;
        END
    END IN6
    PIN IN5
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.86 1.39 3.14 1.76 ;
        END
    END IN5
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.10 1.39 2.38 1.81 ;
        END
    END IN4
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.39 1.62 1.81 ;
        END
    END IN3
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 7.60 3.48 ;
        RECT  7.12 2.88 7.42 3.48 ;
        RECT  7.06 1.84 7.34 2.44 ;
        RECT  7.12 1.84 7.28 3.48 ;
        RECT  6.02 1.84 6.30 2.44 ;
        RECT  6.08 1.84 6.24 3.48 ;
        RECT  3.58 1.92 3.86 2.20 ;
        RECT  3.64 1.92 3.80 3.48 ;
        RECT  1.14 2.02 1.42 2.30 ;
        RECT  1.20 2.02 1.36 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 7.60 0.28 ;
        RECT  7.12 -0.28 7.42 0.32 ;
        RECT  7.06 0.64 7.34 1.24 ;
        RECT  7.12 -0.28 7.28 1.24 ;
        RECT  6.02 0.64 6.30 1.24 ;
        RECT  6.08 -0.28 6.24 1.24 ;
        RECT  4.46 0.63 4.74 0.91 ;
        RECT  4.52 -0.28 4.68 0.91 ;
        RECT  3.42 0.63 3.70 0.91 ;
        RECT  3.48 -0.28 3.64 0.91 ;
        RECT  2.28 0.63 2.56 0.91 ;
        RECT  2.34 -0.28 2.50 0.91 ;
        RECT  1.14 0.63 1.42 0.91 ;
        RECT  1.20 -0.28 1.36 0.91 ;
        RECT  0.10 0.63 0.38 0.91 ;
        RECT  0.16 -0.28 0.32 0.91 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.54 0.63 0.90 0.91 ;
        RECT  0.54 0.63 0.70 2.18 ;
        RECT  0.24 2.02 0.70 2.18 ;
        RECT  0.24 2.02 0.52 2.30 ;
        RECT  0.24 2.02 0.40 2.76 ;
        RECT  0.10 2.48 0.40 2.76 ;
        RECT  1.66 0.63 1.94 0.91 ;
        RECT  1.78 0.63 1.94 2.18 ;
        RECT  1.78 2.02 2.32 2.18 ;
        RECT  2.04 2.02 2.32 2.30 ;
        RECT  2.16 2.02 2.32 2.70 ;
        RECT  2.16 2.42 2.46 2.70 ;
        RECT  2.90 0.63 3.18 0.91 ;
        RECT  2.90 0.63 3.06 1.23 ;
        RECT  2.54 1.07 3.98 1.23 ;
        RECT  3.82 1.07 3.98 1.74 ;
        RECT  3.82 1.46 4.10 1.74 ;
        RECT  2.54 1.07 2.70 2.20 ;
        RECT  2.54 1.92 2.96 2.20 ;
        RECT  3.94 0.63 4.30 0.91 ;
        RECT  4.98 0.63 5.26 0.91 ;
        RECT  4.14 0.63 4.30 1.23 ;
        RECT  4.14 1.07 5.14 1.23 ;
        RECT  4.98 1.40 5.42 1.68 ;
        RECT  4.98 0.63 5.14 2.20 ;
        RECT  4.86 1.92 5.14 2.20 ;
        RECT  5.46 0.70 5.74 1.24 ;
        RECT  5.58 1.46 6.48 1.62 ;
        RECT  6.20 1.40 6.48 1.68 ;
        RECT  5.58 0.70 5.74 2.38 ;
        RECT  5.46 1.84 5.74 2.38 ;
    END
END OR23AND3SP4V1_0

MACRO OR23AND3SP2V1_0
    CLASS CORE ;
    FOREIGN OR23AND3SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 12.90  LAYER ME1  ;
        ANTENNADIFFAREA 5.81  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.44  LAYER ME1  ;
        ANTENNAMAXAREACAR 29.22  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.54 1.84 7.08 2.00 ;
        RECT  6.92 1.08 7.08 2.00 ;
        RECT  6.54 1.08 7.08 1.24 ;
        RECT  6.54 1.84 6.82 2.44 ;
        RECT  6.54 0.64 6.82 1.24 ;
        END
    END OUT
    PIN IN6
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.30 1.39 3.62 1.76 ;
        END
    END IN6
    PIN IN5
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.86 1.39 3.14 1.76 ;
        END
    END IN5
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.10 1.39 2.38 1.81 ;
        END
    END IN4
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.39 1.62 1.81 ;
        END
    END IN3
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 7.20 3.48 ;
        RECT  6.74 2.88 7.02 3.48 ;
        RECT  6.02 1.84 6.30 2.44 ;
        RECT  6.08 1.84 6.24 3.48 ;
        RECT  3.58 1.92 3.86 2.20 ;
        RECT  3.64 1.92 3.80 3.48 ;
        RECT  1.14 2.02 1.42 2.30 ;
        RECT  1.20 2.02 1.36 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 7.20 0.28 ;
        RECT  6.74 -0.28 7.02 0.32 ;
        RECT  6.02 0.64 6.30 1.24 ;
        RECT  6.08 -0.28 6.24 1.24 ;
        RECT  4.46 0.63 4.74 0.91 ;
        RECT  4.52 -0.28 4.68 0.91 ;
        RECT  3.42 0.63 3.70 0.91 ;
        RECT  3.48 -0.28 3.64 0.91 ;
        RECT  2.28 0.63 2.56 0.91 ;
        RECT  2.34 -0.28 2.50 0.91 ;
        RECT  1.14 0.63 1.42 0.91 ;
        RECT  1.20 -0.28 1.36 0.91 ;
        RECT  0.10 0.63 0.38 0.91 ;
        RECT  0.16 -0.28 0.32 0.91 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.54 0.63 0.90 0.91 ;
        RECT  0.54 0.63 0.70 2.18 ;
        RECT  0.24 2.02 0.70 2.18 ;
        RECT  0.24 2.02 0.52 2.30 ;
        RECT  0.24 2.02 0.40 2.76 ;
        RECT  0.10 2.48 0.40 2.76 ;
        RECT  1.66 0.63 1.94 0.91 ;
        RECT  1.78 0.63 1.94 2.18 ;
        RECT  1.78 2.02 2.32 2.18 ;
        RECT  2.04 2.02 2.32 2.30 ;
        RECT  2.16 2.02 2.32 2.70 ;
        RECT  2.16 2.42 2.46 2.70 ;
        RECT  2.90 0.63 3.18 0.91 ;
        RECT  2.90 0.63 3.06 1.23 ;
        RECT  2.54 1.07 3.98 1.23 ;
        RECT  3.82 1.07 3.98 1.74 ;
        RECT  3.82 1.46 4.10 1.74 ;
        RECT  2.54 1.07 2.70 2.20 ;
        RECT  2.54 1.92 2.96 2.20 ;
        RECT  3.94 0.63 4.30 0.91 ;
        RECT  4.96 0.63 5.26 0.91 ;
        RECT  4.14 0.63 4.30 1.23 ;
        RECT  4.14 1.07 5.12 1.23 ;
        RECT  4.96 1.40 5.40 1.68 ;
        RECT  4.96 0.63 5.12 2.20 ;
        RECT  4.86 1.92 5.14 2.20 ;
        RECT  5.46 0.84 5.76 1.24 ;
        RECT  5.60 1.46 6.40 1.62 ;
        RECT  6.12 1.40 6.40 1.68 ;
        RECT  5.60 0.84 5.76 2.24 ;
        RECT  5.46 1.84 5.76 2.24 ;
    END
END OR23AND3SP2V1_0

MACRO OR23AND3SP1V1_0
    CLASS CORE ;
    FOREIGN OR23AND3SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 9.59  LAYER ME1  ;
        ANTENNADIFFAREA 4.14  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.23  LAYER ME1  ;
        ANTENNAMAXAREACAR 41.62  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.92 0.63 5.26 0.91 ;
        RECT  4.90 1.84 5.18 2.20 ;
        RECT  4.92 0.63 5.08 2.20 ;
        RECT  4.14 1.07 5.08 1.23 ;
        RECT  4.14 0.63 4.30 1.23 ;
        RECT  3.94 0.63 4.30 0.91 ;
        END
    END OUT
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN5
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.86 1.39 3.14 1.76 ;
        END
    END IN5
    PIN IN6
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.30 1.39 3.62 1.76 ;
        END
    END IN6
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.10 1.39 2.38 1.81 ;
        END
    END IN4
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.39 1.62 1.81 ;
        END
    END IN3
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 5.60 0.28 ;
        RECT  5.14 -0.28 5.42 0.32 ;
        RECT  4.46 0.63 4.74 0.91 ;
        RECT  4.52 -0.28 4.68 0.91 ;
        RECT  3.42 0.63 3.70 0.91 ;
        RECT  3.48 -0.28 3.64 0.91 ;
        RECT  2.28 0.63 2.56 0.91 ;
        RECT  2.34 -0.28 2.50 0.91 ;
        RECT  1.14 0.63 1.42 0.91 ;
        RECT  1.20 -0.28 1.36 0.91 ;
        RECT  0.10 0.63 0.38 0.91 ;
        RECT  0.16 -0.28 0.32 0.91 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 5.60 3.48 ;
        RECT  5.14 2.88 5.42 3.48 ;
        RECT  3.62 1.92 3.90 2.20 ;
        RECT  3.68 1.92 3.84 3.48 ;
        RECT  1.14 2.02 1.42 2.30 ;
        RECT  1.20 2.02 1.36 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.54 0.63 0.90 0.91 ;
        RECT  0.54 0.63 0.70 2.18 ;
        RECT  0.24 2.02 0.70 2.18 ;
        RECT  0.24 2.02 0.52 2.30 ;
        RECT  0.24 2.02 0.40 2.76 ;
        RECT  0.10 2.48 0.40 2.76 ;
        RECT  1.66 0.63 1.94 0.91 ;
        RECT  1.78 0.63 1.94 2.18 ;
        RECT  1.78 2.02 2.32 2.18 ;
        RECT  2.04 2.02 2.32 2.30 ;
        RECT  2.16 2.02 2.32 2.70 ;
        RECT  2.16 2.42 2.46 2.70 ;
        RECT  2.90 0.63 3.18 0.91 ;
        RECT  2.90 0.63 3.06 1.23 ;
        RECT  2.54 1.07 3.98 1.23 ;
        RECT  3.82 1.07 3.98 1.74 ;
        RECT  3.82 1.46 4.10 1.74 ;
        RECT  2.54 1.07 2.70 2.20 ;
        RECT  2.54 1.92 2.96 2.20 ;
    END
END OR23AND3SP1V1_0

MACRO OR22NAND2SP8V1_0
    CLASS CORE ;
    FOREIGN OR22NAND2SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 11.33  LAYER ME1  ;
        ANTENNADIFFAREA 6.08  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.71  LAYER ME1  ;
        ANTENNAMAXAREACAR 15.95  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.90 1.98 5.18 2.58 ;
        RECT  4.82 0.61 5.10 1.21 ;
        RECT  4.90 0.61 5.06 2.58 ;
        RECT  3.88 1.52 5.06 1.68 ;
        RECT  3.88 1.46 4.32 1.74 ;
        RECT  3.86 1.98 4.14 2.58 ;
        RECT  3.78 0.61 4.06 1.21 ;
        RECT  3.88 0.61 4.04 2.58 ;
        END
    END OUT
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.10 1.47 2.38 1.84 ;
        END
    END IN4
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.36 1.62 1.81 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 6.00 0.28 ;
        RECT  5.40 -0.28 5.82 0.32 ;
        RECT  5.34 0.61 5.62 1.21 ;
        RECT  5.40 -0.28 5.56 1.21 ;
        RECT  4.30 0.61 4.58 1.21 ;
        RECT  4.36 -0.28 4.52 1.21 ;
        RECT  3.26 0.61 3.54 1.21 ;
        RECT  3.32 -0.28 3.48 1.21 ;
        RECT  2.18 0.61 2.46 0.89 ;
        RECT  2.24 -0.28 2.40 0.89 ;
        RECT  1.14 0.61 1.42 0.89 ;
        RECT  1.20 -0.28 1.36 0.89 ;
        RECT  0.10 0.61 0.38 0.89 ;
        RECT  0.16 -0.28 0.32 0.89 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 6.00 3.48 ;
        RECT  5.48 2.88 5.82 3.48 ;
        RECT  5.42 1.98 5.70 2.58 ;
        RECT  5.48 1.98 5.64 3.48 ;
        RECT  4.38 1.98 4.66 2.58 ;
        RECT  4.44 1.98 4.60 3.48 ;
        RECT  3.34 1.98 3.62 2.58 ;
        RECT  3.40 1.98 3.56 3.48 ;
        RECT  1.08 2.02 1.36 2.30 ;
        RECT  1.14 2.02 1.30 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.54 0.61 0.90 0.89 ;
        RECT  0.54 0.61 0.70 2.18 ;
        RECT  0.22 2.02 0.70 2.18 ;
        RECT  0.22 2.02 0.52 2.30 ;
        RECT  0.22 2.02 0.38 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  1.66 0.61 1.94 0.89 ;
        RECT  1.78 1.05 2.74 1.21 ;
        RECT  2.46 1.05 2.74 1.33 ;
        RECT  1.78 0.61 1.94 2.30 ;
        RECT  1.78 2.02 2.20 2.30 ;
        RECT  2.70 0.61 3.06 0.89 ;
        RECT  2.90 1.52 3.72 1.68 ;
        RECT  3.44 1.46 3.72 1.74 ;
        RECT  2.90 0.61 3.06 2.18 ;
        RECT  2.40 2.02 3.06 2.18 ;
        RECT  2.40 2.02 2.68 2.30 ;
    END
END OR22NAND2SP8V1_0

MACRO OR22NAND2SP4V1_0
    CLASS CORE ;
    FOREIGN OR22NAND2SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.36 1.62 1.81 ;
        END
    END IN3
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.10 1.47 2.38 1.84 ;
        END
    END IN4
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.39 0.38 1.81 ;
        END
    END IN1
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 8.98  LAYER ME1  ;
        ANTENNADIFFAREA 4.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.42  LAYER ME1  ;
        ANTENNAMAXAREACAR 21.26  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.88 1.46 4.32 1.74 ;
        RECT  3.86 1.98 4.14 2.58 ;
        RECT  3.78 0.61 4.06 1.21 ;
        RECT  3.88 0.61 4.04 2.58 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.80 3.48 ;
        RECT  4.38 1.98 4.66 2.58 ;
        RECT  4.34 2.88 4.62 3.48 ;
        RECT  4.44 1.98 4.60 3.48 ;
        RECT  3.34 1.98 3.62 2.58 ;
        RECT  3.40 1.98 3.56 3.48 ;
        RECT  1.08 2.02 1.36 2.30 ;
        RECT  1.14 2.02 1.30 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.80 0.28 ;
        RECT  4.34 -0.28 4.62 0.32 ;
        RECT  4.30 0.61 4.58 1.21 ;
        RECT  4.36 -0.28 4.52 1.21 ;
        RECT  3.26 0.61 3.54 1.21 ;
        RECT  3.32 -0.28 3.48 1.21 ;
        RECT  2.18 0.61 2.46 0.89 ;
        RECT  2.24 -0.28 2.40 0.89 ;
        RECT  1.14 0.61 1.42 0.89 ;
        RECT  1.20 -0.28 1.36 0.89 ;
        RECT  0.10 0.61 0.38 0.89 ;
        RECT  0.16 -0.28 0.32 0.89 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.54 0.61 0.90 0.89 ;
        RECT  0.54 0.61 0.70 2.18 ;
        RECT  0.22 2.02 0.70 2.18 ;
        RECT  0.22 2.02 0.52 2.30 ;
        RECT  0.22 2.02 0.38 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  1.66 0.61 1.94 0.89 ;
        RECT  1.78 1.05 2.74 1.21 ;
        RECT  2.46 1.05 2.74 1.33 ;
        RECT  1.78 0.61 1.94 2.30 ;
        RECT  1.78 2.02 2.20 2.30 ;
        RECT  2.70 0.61 3.06 0.89 ;
        RECT  2.90 1.52 3.72 1.68 ;
        RECT  3.44 1.46 3.72 1.74 ;
        RECT  2.90 0.61 3.06 2.18 ;
        RECT  2.40 2.02 3.06 2.18 ;
        RECT  2.40 2.02 2.68 2.30 ;
    END
END OR22NAND2SP4V1_0

MACRO OR22NAND2SP2V1_0
    CLASS CORE ;
    FOREIGN OR22NAND2SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 8.10  LAYER ME1  ;
        ANTENNADIFFAREA 3.76  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.28  LAYER ME1  ;
        ANTENNAMAXAREACAR 29.10  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.88 1.46 4.32 1.74 ;
        RECT  3.86 1.98 4.14 2.58 ;
        RECT  3.78 0.61 4.06 1.21 ;
        RECT  3.88 0.61 4.04 2.58 ;
        END
    END OUT
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.10 1.47 2.38 1.84 ;
        END
    END IN4
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.36 1.62 1.81 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.40 0.28 ;
        RECT  3.94 -0.28 4.22 0.32 ;
        RECT  3.26 0.61 3.54 1.21 ;
        RECT  3.32 -0.28 3.48 1.21 ;
        RECT  2.18 0.61 2.46 0.89 ;
        RECT  2.24 -0.28 2.40 0.89 ;
        RECT  1.14 0.61 1.42 0.89 ;
        RECT  1.20 -0.28 1.36 0.89 ;
        RECT  0.10 0.61 0.38 0.89 ;
        RECT  0.16 -0.28 0.32 0.89 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.40 3.48 ;
        RECT  3.94 2.88 4.22 3.48 ;
        RECT  3.34 1.98 3.62 2.58 ;
        RECT  3.40 1.98 3.56 3.48 ;
        RECT  1.08 2.02 1.36 2.30 ;
        RECT  1.14 2.02 1.30 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.54 0.61 0.90 0.89 ;
        RECT  0.54 0.61 0.70 2.18 ;
        RECT  0.22 2.02 0.70 2.18 ;
        RECT  0.22 2.02 0.52 2.30 ;
        RECT  0.22 2.02 0.38 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  1.66 0.61 1.94 0.89 ;
        RECT  1.78 1.05 2.74 1.21 ;
        RECT  2.46 1.05 2.74 1.33 ;
        RECT  1.78 0.61 1.94 2.30 ;
        RECT  1.78 2.02 2.20 2.30 ;
        RECT  2.70 0.61 3.06 0.89 ;
        RECT  2.90 1.52 3.72 1.68 ;
        RECT  3.44 1.46 3.72 1.74 ;
        RECT  2.90 0.61 3.06 2.18 ;
        RECT  2.40 2.02 3.06 2.18 ;
        RECT  2.40 2.02 2.68 2.30 ;
    END
END OR22NAND2SP2V1_0

MACRO OR22NAND2SP1V1_0
    CLASS CORE ;
    FOREIGN OR22NAND2SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 7.43  LAYER ME1  ;
        ANTENNADIFFAREA 3.31  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        ANTENNAMAXAREACAR 36.86  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.88 1.46 4.32 1.74 ;
        RECT  3.82 2.02 4.10 2.30 ;
        RECT  3.88 0.61 4.04 2.30 ;
        RECT  3.74 0.61 4.04 0.89 ;
        END
    END OUT
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.36 1.62 1.81 ;
        END
    END IN3
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.10 1.47 2.38 1.84 ;
        END
    END IN4
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.40 3.48 ;
        RECT  3.94 2.88 4.22 3.48 ;
        RECT  3.30 2.02 3.58 2.30 ;
        RECT  3.36 2.02 3.52 3.48 ;
        RECT  1.08 2.02 1.36 2.30 ;
        RECT  1.14 2.02 1.30 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.40 0.28 ;
        RECT  3.94 -0.28 4.22 0.32 ;
        RECT  3.22 0.61 3.50 0.89 ;
        RECT  3.28 -0.28 3.44 0.89 ;
        RECT  2.18 0.61 2.46 0.89 ;
        RECT  2.24 -0.28 2.40 0.89 ;
        RECT  1.14 0.61 1.42 0.89 ;
        RECT  1.20 -0.28 1.36 0.89 ;
        RECT  0.10 0.61 0.38 0.89 ;
        RECT  0.16 -0.28 0.32 0.89 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.54 0.61 0.90 0.89 ;
        RECT  0.54 0.61 0.70 2.18 ;
        RECT  0.22 2.02 0.70 2.18 ;
        RECT  0.22 2.02 0.52 2.30 ;
        RECT  0.22 2.02 0.38 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  1.66 0.61 1.94 0.89 ;
        RECT  1.78 1.05 2.74 1.21 ;
        RECT  2.46 1.05 2.74 1.33 ;
        RECT  1.78 0.61 1.94 2.30 ;
        RECT  1.78 2.02 2.20 2.30 ;
        RECT  2.70 0.61 3.06 0.89 ;
        RECT  2.90 1.52 3.72 1.68 ;
        RECT  3.44 1.46 3.72 1.74 ;
        RECT  2.90 0.61 3.06 2.18 ;
        RECT  2.40 2.02 3.06 2.18 ;
        RECT  2.40 2.02 2.68 2.30 ;
    END
END OR22NAND2SP1V1_0

MACRO OR22AND2SP8V1_0
    CLASS CORE ;
    FOREIGN OR22AND2SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 13.92  LAYER ME1  ;
        ANTENNADIFFAREA 7.97  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER ME1  ;
        ANTENNAMAXAREACAR 12.09  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.16 1.92 6.44 2.20 ;
        RECT  6.16 1.46 6.32 2.20 ;
        RECT  5.95 0.63 6.23 1.23 ;
        RECT  6.01 0.63 6.17 1.62 ;
        RECT  3.02 1.46 6.32 1.62 ;
        RECT  5.12 1.92 5.40 2.20 ;
        RECT  5.18 1.46 5.34 2.20 ;
        RECT  4.91 0.63 5.19 1.23 ;
        RECT  4.97 0.63 5.13 1.62 ;
        RECT  3.87 0.63 4.15 1.23 ;
        RECT  3.93 0.63 4.09 1.62 ;
        RECT  3.26 1.46 3.54 1.74 ;
        RECT  3.02 0.69 3.18 1.62 ;
        RECT  2.83 0.69 3.18 0.97 ;
        END
    END OUT
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.10 1.43 2.38 1.84 ;
        END
    END IN4
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.39 1.62 1.81 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 7.20 0.28 ;
        RECT  6.58 -0.28 7.02 0.32 ;
        RECT  6.47 0.63 6.75 1.23 ;
        RECT  6.58 -0.28 6.74 1.23 ;
        RECT  5.43 0.63 5.71 1.23 ;
        RECT  5.49 -0.28 5.65 1.23 ;
        RECT  4.39 0.63 4.67 1.23 ;
        RECT  4.45 -0.28 4.61 1.23 ;
        RECT  3.35 0.63 3.63 1.23 ;
        RECT  3.41 -0.28 3.57 1.23 ;
        RECT  2.31 0.63 2.59 0.91 ;
        RECT  2.37 -0.28 2.53 0.91 ;
        RECT  1.23 0.63 1.51 0.91 ;
        RECT  1.29 -0.28 1.45 0.91 ;
        RECT  0.19 0.63 0.47 0.91 ;
        RECT  0.25 -0.28 0.41 0.91 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 7.20 3.48 ;
        RECT  6.74 2.88 7.02 3.48 ;
        RECT  4.08 2.24 4.36 2.52 ;
        RECT  4.14 2.24 4.30 3.48 ;
        RECT  3.04 2.24 3.32 2.52 ;
        RECT  3.10 2.24 3.26 3.48 ;
        RECT  1.14 2.10 1.42 2.38 ;
        RECT  1.20 2.10 1.36 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.65 0.63 0.99 0.91 ;
        RECT  0.65 0.63 0.81 1.23 ;
        RECT  0.54 1.07 0.70 2.38 ;
        RECT  0.22 2.10 0.70 2.38 ;
        RECT  0.22 2.10 0.38 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  1.75 0.63 2.03 0.91 ;
        RECT  1.78 1.07 2.70 1.23 ;
        RECT  2.54 1.07 2.70 1.67 ;
        RECT  2.54 1.39 2.86 1.67 ;
        RECT  1.78 0.63 1.94 2.26 ;
        RECT  1.78 2.10 2.32 2.26 ;
        RECT  2.04 2.10 2.32 2.38 ;
        RECT  2.52 1.92 4.88 2.08 ;
        RECT  4.60 1.92 4.88 2.52 ;
        RECT  5.64 1.92 5.92 2.52 ;
        RECT  2.52 1.92 2.80 2.52 ;
        RECT  3.56 1.92 3.84 2.52 ;
        RECT  6.68 1.92 6.96 2.52 ;
        RECT  4.60 2.36 6.96 2.52 ;
    END
END OR22AND2SP8V1_0

MACRO OR22AND2SP4V1_0
    CLASS CORE ;
    FOREIGN OR22AND2SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 9.65  LAYER ME1  ;
        ANTENNADIFFAREA 5.41  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.58  LAYER ME1  ;
        ANTENNAMAXAREACAR 16.75  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.08 1.92 4.36 2.20 ;
        RECT  4.08 1.46 4.24 2.20 ;
        RECT  3.87 0.63 4.15 1.23 ;
        RECT  3.93 0.63 4.09 1.62 ;
        RECT  3.02 1.46 4.24 1.62 ;
        RECT  3.26 1.46 3.54 1.74 ;
        RECT  3.02 0.70 3.18 1.62 ;
        RECT  2.83 0.70 3.18 0.97 ;
        END
    END OUT
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.10 1.43 2.38 1.84 ;
        END
    END IN4
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.39 1.62 1.81 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 5.20 0.28 ;
        RECT  4.74 -0.28 5.02 0.32 ;
        RECT  4.39 0.63 4.67 1.23 ;
        RECT  4.42 -0.28 4.58 1.23 ;
        RECT  3.35 0.63 3.63 1.23 ;
        RECT  3.41 -0.28 3.57 1.23 ;
        RECT  2.31 0.63 2.59 0.91 ;
        RECT  2.37 -0.28 2.53 0.91 ;
        RECT  1.23 0.63 1.51 0.91 ;
        RECT  1.29 -0.28 1.45 0.91 ;
        RECT  0.19 0.63 0.47 0.91 ;
        RECT  0.25 -0.28 0.41 0.91 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 5.20 3.48 ;
        RECT  4.74 2.88 5.02 3.48 ;
        RECT  3.04 2.24 3.32 2.52 ;
        RECT  3.10 2.24 3.26 3.48 ;
        RECT  1.14 2.10 1.42 2.38 ;
        RECT  1.20 2.10 1.36 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.65 0.63 0.99 0.91 ;
        RECT  0.65 0.63 0.81 1.23 ;
        RECT  0.54 1.07 0.70 2.38 ;
        RECT  0.22 2.10 0.70 2.38 ;
        RECT  0.22 2.10 0.38 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  1.75 0.63 2.03 0.91 ;
        RECT  1.78 1.07 2.70 1.23 ;
        RECT  2.54 1.07 2.70 1.71 ;
        RECT  2.54 1.43 2.86 1.71 ;
        RECT  1.78 0.63 1.94 2.26 ;
        RECT  1.78 2.10 2.32 2.26 ;
        RECT  2.04 2.10 2.32 2.38 ;
        RECT  2.52 1.92 3.84 2.08 ;
        RECT  3.56 1.92 3.84 2.52 ;
        RECT  2.52 1.92 2.80 2.52 ;
        RECT  4.60 1.92 4.88 2.52 ;
        RECT  3.56 2.36 4.88 2.52 ;
    END
END OR22AND2SP4V1_0

MACRO OR22AND2SP2V1_0
    CLASS CORE ;
    FOREIGN OR22AND2SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 6.68  LAYER ME1  ;
        ANTENNADIFFAREA 3.74  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.29  LAYER ME1  ;
        ANTENNAMAXAREACAR 23.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.38 1.92 3.70 2.52 ;
        RECT  3.38 1.46 3.54 2.52 ;
        RECT  3.26 1.46 3.54 1.74 ;
        RECT  3.02 1.46 3.54 1.62 ;
        RECT  3.02 0.69 3.18 1.62 ;
        RECT  2.83 0.69 3.18 0.97 ;
        END
    END OUT
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.10 1.43 2.38 1.84 ;
        END
    END IN4
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.39 1.62 1.81 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.00 0.28 ;
        RECT  3.41 -0.28 3.82 0.32 ;
        RECT  3.35 0.63 3.63 1.23 ;
        RECT  3.41 -0.28 3.57 1.23 ;
        RECT  2.31 0.63 2.59 0.91 ;
        RECT  2.37 -0.28 2.53 0.91 ;
        RECT  1.23 0.63 1.51 0.91 ;
        RECT  1.29 -0.28 1.45 0.91 ;
        RECT  0.19 0.63 0.47 0.91 ;
        RECT  0.25 -0.28 0.41 0.91 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.00 3.48 ;
        RECT  3.54 2.88 3.82 3.48 ;
        RECT  2.52 1.92 2.80 2.52 ;
        RECT  2.58 1.92 2.74 3.48 ;
        RECT  1.14 2.10 1.42 2.38 ;
        RECT  1.20 2.10 1.36 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.65 0.63 0.99 0.91 ;
        RECT  0.65 0.63 0.81 1.23 ;
        RECT  0.54 1.07 0.70 2.38 ;
        RECT  0.22 2.10 0.70 2.38 ;
        RECT  0.22 2.10 0.38 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  1.75 0.63 2.03 0.91 ;
        RECT  1.78 1.07 2.70 1.23 ;
        RECT  2.54 1.07 2.70 1.66 ;
        RECT  2.54 1.38 2.86 1.66 ;
        RECT  1.78 0.63 1.94 2.26 ;
        RECT  1.78 2.10 2.32 2.26 ;
        RECT  2.04 2.10 2.32 2.38 ;
    END
END OR22AND2SP2V1_0

MACRO OR22AND2SP1V1_0
    CLASS CORE ;
    FOREIGN OR22AND2SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 6.47  LAYER ME1  ;
        ANTENNADIFFAREA 3.08  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        ANTENNAMAXAREACAR 48.11  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.38 2.10 3.70 2.38 ;
        RECT  3.38 1.46 3.54 2.38 ;
        RECT  3.26 1.46 3.54 1.74 ;
        RECT  2.99 1.46 3.54 1.62 ;
        RECT  2.99 0.63 3.15 1.62 ;
        RECT  2.79 0.63 3.15 0.91 ;
        END
    END OUT
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.39 1.62 1.81 ;
        END
    END IN3
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.10 1.43 2.38 1.85 ;
        END
    END IN4
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.00 0.28 ;
        RECT  3.38 -0.28 3.82 0.32 ;
        RECT  3.31 0.63 3.59 0.91 ;
        RECT  3.38 -0.28 3.54 0.91 ;
        RECT  2.27 0.63 2.55 0.91 ;
        RECT  2.33 -0.28 2.49 0.91 ;
        RECT  1.23 0.63 1.51 0.91 ;
        RECT  1.29 -0.28 1.45 0.91 ;
        RECT  0.19 0.63 0.47 0.91 ;
        RECT  0.25 -0.28 0.41 0.91 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.00 3.48 ;
        RECT  3.54 2.88 3.82 3.48 ;
        RECT  2.52 2.10 2.80 2.38 ;
        RECT  2.58 2.10 2.74 3.48 ;
        RECT  1.14 2.10 1.42 2.38 ;
        RECT  1.20 2.10 1.36 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.65 0.63 0.99 0.91 ;
        RECT  0.65 0.63 0.81 1.23 ;
        RECT  0.54 1.07 0.70 2.38 ;
        RECT  0.22 2.10 0.70 2.38 ;
        RECT  0.22 2.10 0.38 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  1.75 0.63 2.03 0.91 ;
        RECT  1.78 1.07 2.83 1.23 ;
        RECT  2.55 1.07 2.83 1.35 ;
        RECT  1.78 0.63 1.94 2.26 ;
        RECT  1.78 2.10 2.32 2.26 ;
        RECT  2.04 2.10 2.32 2.38 ;
    END
END OR22AND2SP1V1_0

MACRO NOR8SP8V1_0
    CLASS CORE ;
    FOREIGN NOR8SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN8
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.10 1.39 8.42 1.81 ;
        END
    END IN8
    PIN IN7
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.66 1.40 7.94 1.81 ;
        END
    END IN7
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 16.13  LAYER ME1  ;
        ANTENNADIFFAREA 8.68  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.91  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.69  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.18 1.90 5.46 2.50 ;
        RECT  5.18 0.63 5.46 1.23 ;
        RECT  5.18 0.63 5.34 2.50 ;
        RECT  4.26 1.52 5.34 1.68 ;
        RECT  4.14 1.90 4.42 2.50 ;
        RECT  4.26 0.63 4.42 2.50 ;
        RECT  4.14 0.63 4.42 1.23 ;
        END
    END OUT
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.39 1.62 1.81 ;
        END
    END IN3
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.10 1.07 2.52 1.35 ;
        END
    END IN4
    PIN IN5
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.06 1.39 6.34 1.81 ;
        END
    END IN5
    PIN IN6
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.90 1.40 7.18 1.81 ;
        END
    END IN6
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 8.80 0.28 ;
        RECT  8.34 -0.28 8.62 0.32 ;
        RECT  7.86 0.63 8.14 0.91 ;
        RECT  7.92 -0.28 8.08 0.91 ;
        RECT  6.82 0.63 7.10 0.91 ;
        RECT  6.89 -0.28 7.05 0.91 ;
        RECT  5.70 0.63 5.98 1.23 ;
        RECT  5.76 -0.28 5.92 1.23 ;
        RECT  4.66 0.63 4.94 1.23 ;
        RECT  4.72 -0.28 4.88 1.23 ;
        RECT  3.58 0.53 3.86 1.23 ;
        RECT  3.64 -0.28 3.80 1.23 ;
        RECT  2.18 0.63 2.46 0.91 ;
        RECT  2.24 -0.28 2.40 0.91 ;
        RECT  1.14 0.63 1.42 0.91 ;
        RECT  1.20 -0.28 1.36 0.91 ;
        RECT  0.10 0.63 0.38 0.91 ;
        RECT  0.16 -0.28 0.32 0.91 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 8.80 3.48 ;
        RECT  8.12 2.88 8.62 3.48 ;
        RECT  8.06 2.10 8.34 2.38 ;
        RECT  8.12 2.10 8.28 3.48 ;
        RECT  5.70 1.96 5.98 2.24 ;
        RECT  5.76 1.96 5.92 3.48 ;
        RECT  4.66 1.90 4.94 2.50 ;
        RECT  4.72 1.90 4.88 3.48 ;
        RECT  3.58 1.90 3.86 2.60 ;
        RECT  3.64 1.90 3.80 3.48 ;
        RECT  2.54 1.90 2.82 2.60 ;
        RECT  2.60 1.90 2.76 3.48 ;
        RECT  0.24 2.08 0.52 2.36 ;
        RECT  0.30 2.08 0.46 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.63 0.90 0.91 ;
        RECT  1.66 0.63 1.94 0.91 ;
        RECT  0.74 0.63 0.90 1.23 ;
        RECT  0.74 1.07 1.94 1.23 ;
        RECT  2.75 1.46 3.03 1.74 ;
        RECT  1.78 1.58 3.03 1.74 ;
        RECT  1.78 0.63 1.94 2.36 ;
        RECT  1.78 2.08 2.18 2.36 ;
        RECT  2.68 0.53 2.96 1.23 ;
        RECT  2.68 1.07 3.35 1.23 ;
        RECT  3.19 1.52 4.00 1.68 ;
        RECT  3.72 1.46 4.00 1.74 ;
        RECT  3.19 1.07 3.35 2.60 ;
        RECT  3.06 1.90 3.35 2.60 ;
        RECT  6.21 0.63 6.58 0.91 ;
        RECT  7.34 0.63 7.62 0.91 ;
        RECT  8.38 0.63 8.66 0.91 ;
        RECT  6.21 0.63 6.37 1.23 ;
        RECT  7.40 0.63 7.56 1.23 ;
        RECT  8.38 0.63 8.54 1.23 ;
        RECT  6.21 1.07 8.54 1.23 ;
        RECT  6.52 1.07 6.68 2.38 ;
        RECT  6.28 2.10 6.68 2.38 ;
        RECT  6.28 2.10 6.44 2.76 ;
        RECT  6.08 2.48 6.44 2.76 ;
    END
END NOR8SP8V1_0

MACRO NOR8SP4V1_0
    CLASS CORE ;
    FOREIGN NOR8SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN6
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.70 1.40 6.14 1.74 ;
        END
    END IN6
    PIN IN5
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.26 1.39 5.54 1.81 ;
        END
    END IN5
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.10 1.07 2.52 1.35 ;
        END
    END IN4
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.39 1.62 1.81 ;
        END
    END IN3
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 13.80  LAYER ME1  ;
        ANTENNADIFFAREA 6.75  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER ME1  ;
        ANTENNAMAXAREACAR 24.37  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.26 1.52 4.68 1.68 ;
        RECT  4.14 1.90 4.42 2.50 ;
        RECT  4.26 0.63 4.42 2.50 ;
        RECT  4.14 0.63 4.42 1.23 ;
        END
    END OUT
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN7
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.62 1.40 7.14 1.73 ;
        END
    END IN7
    PIN IN8
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.30 1.39 7.58 1.81 ;
        END
    END IN8
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 8.00 0.28 ;
        RECT  7.54 -0.28 7.82 0.32 ;
        RECT  6.82 0.63 7.10 0.91 ;
        RECT  6.88 -0.28 7.04 0.91 ;
        RECT  5.78 0.63 6.06 0.91 ;
        RECT  5.85 -0.28 6.01 0.91 ;
        RECT  4.66 0.63 4.94 1.23 ;
        RECT  4.72 -0.28 4.88 1.23 ;
        RECT  3.62 0.63 3.90 1.23 ;
        RECT  3.68 -0.28 3.84 1.23 ;
        RECT  2.18 0.63 2.46 0.91 ;
        RECT  2.24 -0.28 2.40 0.91 ;
        RECT  1.14 0.63 1.42 0.91 ;
        RECT  1.20 -0.28 1.36 0.91 ;
        RECT  0.10 0.63 0.38 0.91 ;
        RECT  0.16 -0.28 0.32 0.91 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 8.00 3.48 ;
        RECT  7.54 2.88 7.82 3.48 ;
        RECT  7.02 2.10 7.30 2.38 ;
        RECT  7.08 2.10 7.24 3.48 ;
        RECT  4.66 1.90 4.94 2.18 ;
        RECT  4.72 1.90 4.88 3.48 ;
        RECT  3.62 1.90 3.90 2.50 ;
        RECT  3.68 1.90 3.84 3.48 ;
        RECT  2.54 1.90 2.82 2.48 ;
        RECT  2.60 1.90 2.76 3.48 ;
        RECT  0.24 2.08 0.52 2.36 ;
        RECT  0.30 2.08 0.46 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.63 0.90 0.91 ;
        RECT  1.66 0.63 1.94 0.91 ;
        RECT  0.74 0.63 0.90 1.23 ;
        RECT  0.74 1.07 1.94 1.23 ;
        RECT  2.75 1.46 3.03 1.74 ;
        RECT  1.78 1.58 3.03 1.74 ;
        RECT  1.78 0.63 1.94 2.36 ;
        RECT  1.78 2.08 2.18 2.36 ;
        RECT  2.68 0.65 2.96 1.23 ;
        RECT  2.68 1.07 3.35 1.23 ;
        RECT  3.19 1.52 4.00 1.68 ;
        RECT  3.72 1.46 4.00 1.74 ;
        RECT  3.19 1.07 3.35 2.30 ;
        RECT  3.06 1.90 3.34 2.48 ;
        RECT  5.17 0.63 5.54 0.91 ;
        RECT  6.30 0.63 6.58 0.91 ;
        RECT  7.34 0.63 7.62 0.91 ;
        RECT  5.17 0.63 5.33 1.23 ;
        RECT  6.36 0.63 6.52 1.23 ;
        RECT  7.34 0.63 7.50 1.23 ;
        RECT  5.17 1.07 7.50 1.23 ;
        RECT  6.30 1.07 6.46 2.26 ;
        RECT  5.24 2.10 6.46 2.26 ;
        RECT  5.24 2.10 5.64 2.38 ;
        RECT  5.24 2.10 5.40 2.76 ;
        RECT  5.04 2.48 5.40 2.76 ;
    END
END NOR8SP4V1_0

MACRO NOR8SP2V1_0
    CLASS CORE ;
    FOREIGN NOR8SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN8
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.82 1.39 7.10 1.81 ;
        END
    END IN8
    PIN IN7
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.10 1.40 6.38 1.81 ;
        END
    END IN7
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 12.36  LAYER ME1  ;
        ANTENNADIFFAREA 5.74  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.34  LAYER ME1  ;
        ANTENNAMAXAREACAR 36.79  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.26 1.52 4.68 1.68 ;
        RECT  4.14 1.90 4.42 2.18 ;
        RECT  4.26 0.63 4.42 2.18 ;
        RECT  4.14 0.63 4.42 1.23 ;
        END
    END OUT
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.39 1.62 1.81 ;
        END
    END IN3
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.10 1.07 2.52 1.35 ;
        END
    END IN4
    PIN IN5
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.86 1.39 5.14 1.81 ;
        END
    END IN5
    PIN IN6
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.30 1.40 5.62 1.81 ;
        END
    END IN6
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 7.20 3.48 ;
        RECT  6.56 2.88 7.02 3.48 ;
        RECT  6.50 2.10 6.78 2.38 ;
        RECT  6.56 2.10 6.72 3.48 ;
        RECT  3.62 1.90 3.90 2.50 ;
        RECT  3.68 1.90 3.84 3.48 ;
        RECT  2.54 1.90 2.82 2.30 ;
        RECT  2.60 1.90 2.76 3.48 ;
        RECT  0.24 2.08 0.52 2.36 ;
        RECT  0.30 2.08 0.46 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 7.20 0.28 ;
        RECT  6.74 -0.28 7.02 0.32 ;
        RECT  6.30 0.63 6.58 0.91 ;
        RECT  6.36 -0.28 6.52 0.91 ;
        RECT  5.26 0.63 5.54 0.91 ;
        RECT  5.33 -0.28 5.49 0.91 ;
        RECT  3.62 0.63 3.90 1.23 ;
        RECT  3.68 -0.28 3.84 1.23 ;
        RECT  2.18 0.63 2.46 0.91 ;
        RECT  2.24 -0.28 2.40 0.91 ;
        RECT  1.14 0.63 1.42 0.91 ;
        RECT  1.20 -0.28 1.36 0.91 ;
        RECT  0.10 0.63 0.38 0.91 ;
        RECT  0.16 -0.28 0.32 0.91 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.63 0.90 0.91 ;
        RECT  1.66 0.63 1.94 0.91 ;
        RECT  0.74 0.63 0.90 1.23 ;
        RECT  0.74 1.07 1.94 1.23 ;
        RECT  2.75 1.46 3.03 1.74 ;
        RECT  1.78 1.58 3.03 1.74 ;
        RECT  1.78 0.63 1.94 2.36 ;
        RECT  1.78 2.08 2.18 2.36 ;
        RECT  2.68 0.83 2.96 1.23 ;
        RECT  2.68 1.07 3.35 1.23 ;
        RECT  3.19 1.52 4.00 1.68 ;
        RECT  3.72 1.46 4.00 1.74 ;
        RECT  3.19 1.07 3.35 2.30 ;
        RECT  3.06 1.90 3.35 2.30 ;
        RECT  4.65 0.63 5.02 0.91 ;
        RECT  5.78 0.63 6.06 0.91 ;
        RECT  6.82 0.63 7.10 0.91 ;
        RECT  4.65 0.63 4.81 1.23 ;
        RECT  5.84 0.63 6.00 1.23 ;
        RECT  6.82 0.63 6.98 1.23 ;
        RECT  4.65 1.07 6.98 1.23 ;
        RECT  5.78 1.07 5.94 2.26 ;
        RECT  4.72 2.10 5.94 2.26 ;
        RECT  4.72 2.10 5.12 2.38 ;
        RECT  4.72 2.10 4.88 2.76 ;
        RECT  4.52 2.48 4.88 2.76 ;
    END
END NOR8SP2V1_0

MACRO NOR8SP1V1_0
    CLASS CORE ;
    FOREIGN NOR8SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN6
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.30 1.39 5.62 1.81 ;
        END
    END IN6
    PIN IN5
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.86 1.39 5.14 1.81 ;
        END
    END IN5
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.10 1.07 2.52 1.35 ;
        END
    END IN4
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.39 1.62 1.81 ;
        END
    END IN3
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 12.43  LAYER ME1  ;
        ANTENNADIFFAREA 5.10  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        ANTENNAMAXAREACAR 61.63  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.19 1.52 4.68 1.68 ;
        RECT  4.13 1.90 4.41 2.18 ;
        RECT  4.10 0.95 4.38 1.23 ;
        RECT  4.19 0.95 4.35 2.18 ;
        END
    END OUT
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN7
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.00 1.39 6.28 1.81 ;
        END
    END IN7
    PIN IN8
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.48 1.39 6.76 1.81 ;
        END
    END IN8
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 7.20 0.28 ;
        RECT  6.74 -0.28 7.02 0.32 ;
        RECT  6.24 0.63 6.52 0.91 ;
        RECT  6.30 -0.28 6.46 0.91 ;
        RECT  5.20 0.63 5.48 0.91 ;
        RECT  5.27 -0.28 5.43 0.91 ;
        RECT  3.58 0.95 3.86 1.23 ;
        RECT  3.64 -0.28 3.80 1.23 ;
        RECT  2.18 0.63 2.46 0.91 ;
        RECT  2.24 -0.28 2.40 0.91 ;
        RECT  1.14 0.63 1.42 0.91 ;
        RECT  1.20 -0.28 1.36 0.91 ;
        RECT  0.10 0.63 0.38 0.91 ;
        RECT  0.16 -0.28 0.32 0.91 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 7.20 3.48 ;
        RECT  6.50 2.88 7.02 3.48 ;
        RECT  6.44 2.29 6.72 2.57 ;
        RECT  6.50 2.29 6.66 3.48 ;
        RECT  3.61 1.90 3.89 2.18 ;
        RECT  3.71 1.90 3.87 3.48 ;
        RECT  2.57 1.90 2.85 2.18 ;
        RECT  2.63 1.90 2.79 3.48 ;
        RECT  0.24 2.08 0.52 2.36 ;
        RECT  0.30 2.08 0.46 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.63 0.90 0.91 ;
        RECT  1.66 0.63 1.94 0.91 ;
        RECT  0.74 0.63 0.90 1.23 ;
        RECT  0.74 1.07 1.94 1.23 ;
        RECT  2.75 1.46 3.03 1.74 ;
        RECT  1.78 1.58 3.03 1.74 ;
        RECT  1.78 0.63 1.94 2.36 ;
        RECT  1.78 2.08 2.18 2.36 ;
        RECT  2.68 0.95 2.96 1.23 ;
        RECT  2.68 1.07 3.35 1.23 ;
        RECT  3.19 1.52 4.03 1.68 ;
        RECT  3.75 1.46 4.03 1.74 ;
        RECT  3.19 1.07 3.35 2.18 ;
        RECT  3.09 1.90 3.37 2.18 ;
        RECT  4.68 0.63 4.96 0.91 ;
        RECT  5.72 0.63 6.00 0.91 ;
        RECT  6.76 0.63 7.04 0.91 ;
        RECT  4.57 0.64 4.73 1.23 ;
        RECT  5.78 0.63 5.94 1.23 ;
        RECT  6.76 0.63 6.92 1.23 ;
        RECT  4.57 1.07 7.08 1.23 ;
        RECT  6.92 1.07 7.08 2.13 ;
        RECT  4.78 1.97 7.08 2.13 ;
        RECT  4.78 1.97 4.94 2.64 ;
        RECT  4.78 2.29 5.06 2.64 ;
        RECT  4.34 2.48 5.06 2.64 ;
        RECT  4.34 2.48 4.62 2.76 ;
    END
END NOR8SP1V1_0

MACRO NOR6SP8V1_0
    CLASS CORE ;
    FOREIGN NOR6SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN6
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.26 1.39 7.54 1.81 ;
        END
    END IN6
    PIN IN5
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.50 1.39 6.90 1.81 ;
        END
    END IN5
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.06 1.39 6.34 1.81 ;
        END
    END IN4
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 14.86  LAYER ME1  ;
        ANTENNADIFFAREA 8.28  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.91  LAYER ME1  ;
        ANTENNAMAXAREACAR 16.30  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.74 1.90 5.02 2.50 ;
        RECT  4.71 0.63 4.99 1.23 ;
        RECT  4.74 0.63 4.90 2.50 ;
        RECT  3.72 1.52 4.90 1.68 ;
        RECT  3.70 1.90 3.98 2.50 ;
        RECT  3.67 0.63 3.95 1.23 ;
        RECT  3.72 0.63 3.88 2.50 ;
        END
    END OUT
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.39 1.62 1.81 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 8.00 3.48 ;
        RECT  7.30 2.88 7.82 3.48 ;
        RECT  7.24 2.10 7.52 2.38 ;
        RECT  7.30 2.10 7.46 3.48 ;
        RECT  5.26 1.90 5.54 2.18 ;
        RECT  5.32 1.90 5.48 3.48 ;
        RECT  4.22 1.90 4.50 2.50 ;
        RECT  4.28 1.90 4.44 3.48 ;
        RECT  3.14 1.90 3.42 2.60 ;
        RECT  3.20 1.90 3.36 3.48 ;
        RECT  2.10 1.90 2.38 2.60 ;
        RECT  2.16 1.90 2.32 3.48 ;
        RECT  0.24 2.08 0.52 2.36 ;
        RECT  0.30 2.08 0.46 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 8.00 0.28 ;
        RECT  7.48 -0.28 7.82 0.32 ;
        RECT  7.42 0.63 7.70 0.91 ;
        RECT  7.48 -0.28 7.64 0.91 ;
        RECT  6.38 0.63 6.66 0.91 ;
        RECT  6.45 -0.28 6.61 0.91 ;
        RECT  5.23 0.63 5.51 1.23 ;
        RECT  5.29 -0.28 5.45 1.23 ;
        RECT  4.19 0.63 4.47 1.23 ;
        RECT  4.25 -0.28 4.41 1.23 ;
        RECT  3.11 0.53 3.39 1.23 ;
        RECT  3.17 -0.28 3.33 1.23 ;
        RECT  1.14 0.63 1.42 0.91 ;
        RECT  1.20 -0.28 1.36 0.91 ;
        RECT  0.10 0.63 0.38 0.91 ;
        RECT  0.16 -0.28 0.32 0.91 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.63 0.90 0.91 ;
        RECT  1.66 0.63 1.94 0.91 ;
        RECT  0.74 0.63 0.90 1.23 ;
        RECT  0.74 1.07 1.94 1.23 ;
        RECT  1.78 1.52 2.56 1.68 ;
        RECT  2.28 1.46 2.56 1.74 ;
        RECT  1.78 0.63 1.94 2.36 ;
        RECT  1.52 2.08 1.94 2.36 ;
        RECT  2.21 0.53 2.49 1.23 ;
        RECT  2.21 1.07 2.88 1.23 ;
        RECT  2.72 1.52 3.56 1.68 ;
        RECT  3.28 1.46 3.56 1.74 ;
        RECT  2.72 1.07 2.88 2.60 ;
        RECT  2.62 1.90 2.90 2.60 ;
        RECT  5.70 0.63 6.14 0.91 ;
        RECT  6.90 0.63 7.18 0.91 ;
        RECT  5.70 0.63 5.86 1.23 ;
        RECT  7.02 0.63 7.18 1.23 ;
        RECT  5.70 1.07 7.18 1.23 ;
        RECT  5.74 1.07 5.90 2.76 ;
        RECT  5.74 2.10 6.24 2.38 ;
        RECT  5.74 2.10 6.00 2.76 ;
        RECT  5.68 2.48 6.00 2.76 ;
    END
END NOR6SP8V1_0

MACRO NOR6SP4V1_0
    CLASS CORE ;
    FOREIGN NOR6SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.39 1.62 1.81 ;
        END
    END IN3
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.86 1.39 5.14 1.81 ;
        END
    END IN4
    PIN IN5
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.64 1.39 5.94 1.81 ;
        END
    END IN5
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 11.92  LAYER ME1  ;
        ANTENNADIFFAREA 6.22  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER ME1  ;
        ANTENNAMAXAREACAR 21.05  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.70 1.90 3.98 2.50 ;
        RECT  3.67 0.63 3.95 1.23 ;
        RECT  3.72 0.63 3.88 2.50 ;
        END
    END OUT
    PIN IN6
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.10 1.39 6.42 1.81 ;
        END
    END IN6
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 6.80 3.48 ;
        RECT  6.26 2.88 6.62 3.48 ;
        RECT  6.20 2.10 6.48 2.38 ;
        RECT  6.26 2.10 6.42 3.48 ;
        RECT  4.22 1.90 4.50 2.18 ;
        RECT  4.28 1.90 4.44 3.48 ;
        RECT  3.18 1.90 3.46 2.50 ;
        RECT  3.24 1.90 3.40 3.48 ;
        RECT  2.10 1.90 2.38 2.48 ;
        RECT  2.16 1.90 2.32 3.48 ;
        RECT  0.24 2.08 0.52 2.36 ;
        RECT  0.30 2.08 0.46 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 6.80 0.28 ;
        RECT  6.38 0.63 6.66 0.91 ;
        RECT  6.34 -0.28 6.62 0.32 ;
        RECT  6.44 -0.28 6.60 0.91 ;
        RECT  5.34 0.63 5.62 0.91 ;
        RECT  5.41 -0.28 5.57 0.91 ;
        RECT  4.19 0.63 4.47 1.23 ;
        RECT  4.25 -0.28 4.41 1.23 ;
        RECT  3.15 0.63 3.43 1.23 ;
        RECT  3.21 -0.28 3.37 1.23 ;
        RECT  1.14 0.63 1.42 0.91 ;
        RECT  1.20 -0.28 1.36 0.91 ;
        RECT  0.10 0.63 0.38 0.91 ;
        RECT  0.16 -0.28 0.32 0.91 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.63 0.90 0.91 ;
        RECT  1.66 0.63 1.94 0.91 ;
        RECT  0.74 0.63 0.90 1.23 ;
        RECT  0.74 1.07 1.94 1.23 ;
        RECT  1.78 1.52 2.56 1.68 ;
        RECT  2.28 1.46 2.56 1.74 ;
        RECT  1.78 0.63 1.94 2.36 ;
        RECT  1.52 2.08 1.94 2.36 ;
        RECT  2.21 0.65 2.49 1.23 ;
        RECT  2.21 1.07 2.88 1.23 ;
        RECT  2.72 1.52 3.56 1.68 ;
        RECT  3.28 1.46 3.56 1.74 ;
        RECT  2.72 1.07 2.88 2.48 ;
        RECT  2.62 1.90 2.90 2.48 ;
        RECT  4.66 0.63 5.10 0.91 ;
        RECT  5.86 0.63 6.14 0.91 ;
        RECT  4.66 0.63 4.82 1.23 ;
        RECT  5.98 0.63 6.14 1.23 ;
        RECT  4.66 1.07 6.14 1.23 ;
        RECT  5.30 1.07 5.46 2.26 ;
        RECT  4.80 2.10 5.46 2.26 ;
        RECT  4.80 2.10 5.20 2.38 ;
        RECT  4.80 2.10 4.96 2.76 ;
        RECT  4.64 2.48 4.96 2.76 ;
    END
END NOR6SP4V1_0

MACRO NOR6SP2V1_0
    CLASS CORE ;
    FOREIGN NOR6SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN6
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.66 1.39 5.94 1.81 ;
        END
    END IN6
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 10.87  LAYER ME1  ;
        ANTENNADIFFAREA 5.34  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.34  LAYER ME1  ;
        ANTENNAMAXAREACAR 32.34  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.70 1.90 3.98 2.18 ;
        RECT  3.67 0.63 3.95 1.23 ;
        RECT  3.72 0.63 3.88 2.18 ;
        END
    END OUT
    PIN IN5
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.90 1.39 5.22 1.81 ;
        END
    END IN5
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.46 1.39 4.74 1.81 ;
        END
    END IN4
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.39 1.62 1.81 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 6.40 0.28 ;
        RECT  5.80 -0.28 6.22 0.32 ;
        RECT  5.74 0.63 6.02 0.91 ;
        RECT  5.80 -0.28 5.96 0.91 ;
        RECT  4.70 0.63 4.98 0.91 ;
        RECT  4.77 -0.28 4.93 0.91 ;
        RECT  3.15 0.63 3.43 1.23 ;
        RECT  3.21 -0.28 3.37 1.23 ;
        RECT  1.14 0.63 1.42 0.91 ;
        RECT  1.20 -0.28 1.36 0.91 ;
        RECT  0.10 0.63 0.38 0.91 ;
        RECT  0.16 -0.28 0.32 0.91 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 6.40 3.48 ;
        RECT  5.94 2.88 6.22 3.48 ;
        RECT  5.56 2.10 5.84 2.38 ;
        RECT  5.62 2.10 5.78 3.48 ;
        RECT  3.18 1.90 3.46 2.50 ;
        RECT  3.24 1.90 3.40 3.48 ;
        RECT  2.10 1.90 2.38 2.30 ;
        RECT  2.16 1.90 2.32 3.48 ;
        RECT  0.24 2.08 0.52 2.36 ;
        RECT  0.30 2.08 0.46 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.63 0.90 0.91 ;
        RECT  1.66 0.63 1.94 0.91 ;
        RECT  0.74 0.63 0.90 1.23 ;
        RECT  0.74 1.07 1.94 1.23 ;
        RECT  1.78 1.52 2.56 1.68 ;
        RECT  2.28 1.46 2.56 1.74 ;
        RECT  1.78 0.63 1.94 2.36 ;
        RECT  1.52 2.08 1.94 2.36 ;
        RECT  2.21 0.83 2.49 1.23 ;
        RECT  2.21 1.07 2.88 1.23 ;
        RECT  2.72 1.52 3.56 1.68 ;
        RECT  3.28 1.46 3.56 1.74 ;
        RECT  2.72 1.07 2.88 2.30 ;
        RECT  2.62 1.90 2.90 2.30 ;
        RECT  4.14 0.63 4.46 0.91 ;
        RECT  5.22 0.63 5.50 0.91 ;
        RECT  5.34 0.63 5.50 1.23 ;
        RECT  4.14 1.07 5.50 1.23 ;
        RECT  4.14 0.63 4.30 2.76 ;
        RECT  4.14 2.10 4.56 2.38 ;
        RECT  4.14 2.10 4.44 2.76 ;
        RECT  4.12 2.48 4.44 2.76 ;
    END
END NOR6SP2V1_0

MACRO NOR6SP1V1_0
    CLASS CORE ;
    FOREIGN NOR6SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 10.71  LAYER ME1  ;
        ANTENNADIFFAREA 4.70  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        ANTENNAMAXAREACAR 53.11  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.66 1.90 3.94 2.18 ;
        RECT  3.63 0.95 3.91 1.23 ;
        RECT  3.72 0.95 3.88 2.18 ;
        END
    END OUT
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.39 1.62 1.81 ;
        END
    END IN3
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.46 1.39 4.74 1.81 ;
        END
    END IN4
    PIN IN5
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.90 1.39 5.22 1.81 ;
        END
    END IN5
    PIN IN6
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.66 1.39 5.94 1.81 ;
        END
    END IN6
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 6.40 3.48 ;
        RECT  5.94 2.88 6.22 3.48 ;
        RECT  5.56 2.10 5.84 2.38 ;
        RECT  5.62 2.10 5.78 3.48 ;
        RECT  3.14 1.90 3.42 2.18 ;
        RECT  3.24 1.90 3.40 3.48 ;
        RECT  2.10 1.90 2.38 2.18 ;
        RECT  2.16 1.90 2.32 3.48 ;
        RECT  0.24 2.08 0.52 2.36 ;
        RECT  0.30 2.08 0.46 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 6.40 0.28 ;
        RECT  5.80 -0.28 6.22 0.32 ;
        RECT  5.74 0.63 6.02 0.91 ;
        RECT  5.80 -0.28 5.96 0.91 ;
        RECT  4.70 0.63 4.98 0.91 ;
        RECT  4.77 -0.28 4.93 0.91 ;
        RECT  3.11 0.95 3.39 1.23 ;
        RECT  3.17 -0.28 3.33 1.23 ;
        RECT  1.14 0.63 1.42 0.91 ;
        RECT  1.20 -0.28 1.36 0.91 ;
        RECT  0.10 0.63 0.38 0.91 ;
        RECT  0.16 -0.28 0.32 0.91 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.63 0.90 0.91 ;
        RECT  1.66 0.63 1.94 0.91 ;
        RECT  0.74 0.63 0.90 1.23 ;
        RECT  0.74 1.07 1.94 1.23 ;
        RECT  1.78 1.52 2.56 1.68 ;
        RECT  2.28 1.46 2.56 1.74 ;
        RECT  1.78 0.63 1.94 2.36 ;
        RECT  1.52 2.08 1.94 2.36 ;
        RECT  2.21 0.95 2.49 1.23 ;
        RECT  2.21 1.07 2.88 1.23 ;
        RECT  2.72 1.52 3.56 1.68 ;
        RECT  3.28 1.46 3.56 1.74 ;
        RECT  2.72 1.07 2.88 2.18 ;
        RECT  2.62 1.90 2.90 2.18 ;
        RECT  4.14 0.63 4.46 0.91 ;
        RECT  5.22 0.63 5.50 0.91 ;
        RECT  5.34 0.63 5.50 1.23 ;
        RECT  4.14 1.07 5.50 1.23 ;
        RECT  4.14 0.63 4.30 2.76 ;
        RECT  4.14 2.10 4.56 2.38 ;
        RECT  4.14 2.10 4.44 2.76 ;
        RECT  4.12 2.48 4.44 2.76 ;
    END
END NOR6SP1V1_0

MACRO NOR5SP8V1_0
    CLASS CORE ;
    FOREIGN NOR5SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 13.67  LAYER ME1  ;
        ANTENNADIFFAREA 7.73  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.91  LAYER ME1  ;
        ANTENNAMAXAREACAR 14.99  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.78 1.90 5.06 2.50 ;
        RECT  4.71 0.63 4.99 1.23 ;
        RECT  4.78 0.63 4.94 2.50 ;
        RECT  3.84 1.52 4.94 1.68 ;
        RECT  3.74 1.90 4.02 2.50 ;
        RECT  3.84 0.63 4.00 2.50 ;
        RECT  3.67 0.63 4.00 1.23 ;
        END
    END OUT
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.39 1.62 1.81 ;
        END
    END IN3
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.66 1.39 5.94 1.81 ;
        END
    END IN4
    PIN IN5
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.82 1.39 7.10 1.81 ;
        END
    END IN5
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 7.20 3.48 ;
        RECT  6.74 2.88 7.02 3.48 ;
        RECT  6.72 1.97 7.00 2.25 ;
        RECT  6.78 1.97 6.94 3.48 ;
        RECT  5.30 2.07 5.58 2.35 ;
        RECT  5.36 2.07 5.52 3.48 ;
        RECT  4.26 1.90 4.54 2.50 ;
        RECT  4.32 1.90 4.48 3.48 ;
        RECT  3.18 1.90 3.46 2.60 ;
        RECT  3.24 1.90 3.40 3.48 ;
        RECT  2.14 1.90 2.42 2.60 ;
        RECT  2.20 1.90 2.36 3.48 ;
        RECT  0.24 2.08 0.52 2.36 ;
        RECT  0.30 2.08 0.46 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 7.20 0.28 ;
        RECT  6.78 0.95 7.06 1.23 ;
        RECT  6.74 -0.28 7.02 0.32 ;
        RECT  6.84 -0.28 7.00 1.23 ;
        RECT  5.74 0.95 6.02 1.23 ;
        RECT  5.80 -0.28 5.96 1.23 ;
        RECT  5.23 0.63 5.51 1.23 ;
        RECT  5.29 -0.28 5.45 1.23 ;
        RECT  4.19 0.63 4.47 1.23 ;
        RECT  4.25 -0.28 4.41 1.23 ;
        RECT  3.11 0.53 3.39 1.23 ;
        RECT  3.17 -0.28 3.33 1.23 ;
        RECT  1.14 0.63 1.42 0.91 ;
        RECT  1.20 -0.28 1.36 0.91 ;
        RECT  0.10 0.63 0.38 0.91 ;
        RECT  0.16 -0.28 0.32 0.91 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.63 0.90 0.91 ;
        RECT  1.66 0.63 1.94 0.91 ;
        RECT  0.74 0.63 0.90 1.23 ;
        RECT  0.74 1.07 1.94 1.23 ;
        RECT  1.78 1.52 2.56 1.68 ;
        RECT  2.28 1.46 2.56 1.74 ;
        RECT  1.78 0.63 1.94 2.36 ;
        RECT  1.52 2.08 1.94 2.36 ;
        RECT  2.21 0.53 2.49 1.23 ;
        RECT  2.21 1.07 2.88 1.23 ;
        RECT  2.72 1.52 3.68 1.68 ;
        RECT  3.40 1.46 3.68 1.74 ;
        RECT  2.72 1.07 2.88 2.60 ;
        RECT  2.66 1.90 2.94 2.60 ;
        RECT  6.22 0.95 6.54 1.23 ;
        RECT  6.22 0.95 6.38 2.13 ;
        RECT  5.82 1.97 6.38 2.13 ;
        RECT  5.82 1.97 6.10 2.25 ;
        RECT  5.88 1.97 6.04 2.76 ;
        RECT  5.68 2.48 6.04 2.76 ;
    END
END NOR5SP8V1_0

MACRO NOR5SP4V1_0
    CLASS CORE ;
    FOREIGN NOR5SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN5
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.66 1.39 5.94 1.81 ;
        END
    END IN5
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.86 1.39 5.14 1.81 ;
        END
    END IN4
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.39 1.62 1.81 ;
        END
    END IN3
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 11.72  LAYER ME1  ;
        ANTENNADIFFAREA 5.80  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER ME1  ;
        ANTENNAMAXAREACAR 20.69  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.86 1.52 4.28 1.68 ;
        RECT  3.74 1.90 4.02 2.50 ;
        RECT  3.86 0.63 4.02 2.50 ;
        RECT  3.67 0.63 4.02 1.23 ;
        END
    END OUT
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 6.40 0.28 ;
        RECT  5.80 -0.28 6.22 0.32 ;
        RECT  5.74 0.95 6.02 1.23 ;
        RECT  5.80 -0.28 5.96 1.23 ;
        RECT  4.70 0.95 4.98 1.23 ;
        RECT  4.76 -0.28 4.92 1.23 ;
        RECT  4.19 0.63 4.47 1.23 ;
        RECT  4.25 -0.28 4.41 1.23 ;
        RECT  3.15 0.63 3.43 1.23 ;
        RECT  3.21 -0.28 3.37 1.23 ;
        RECT  1.14 0.63 1.42 0.91 ;
        RECT  1.20 -0.28 1.36 0.91 ;
        RECT  0.10 0.63 0.38 0.91 ;
        RECT  0.16 -0.28 0.32 0.91 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 6.40 3.48 ;
        RECT  5.74 2.88 6.22 3.48 ;
        RECT  5.68 1.97 5.96 2.25 ;
        RECT  5.74 1.97 5.90 3.48 ;
        RECT  4.26 2.06 4.54 2.34 ;
        RECT  4.32 2.06 4.48 3.48 ;
        RECT  3.21 1.90 3.49 2.50 ;
        RECT  3.27 1.90 3.43 3.48 ;
        RECT  2.14 1.90 2.42 2.48 ;
        RECT  2.20 1.90 2.36 3.48 ;
        RECT  0.24 2.08 0.52 2.36 ;
        RECT  0.30 2.08 0.46 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.63 0.90 0.91 ;
        RECT  1.66 0.63 1.94 0.91 ;
        RECT  0.74 0.63 0.90 1.23 ;
        RECT  0.74 1.07 1.94 1.23 ;
        RECT  1.78 1.52 2.56 1.68 ;
        RECT  2.28 1.46 2.56 1.74 ;
        RECT  1.78 0.63 1.94 2.36 ;
        RECT  1.52 2.08 1.94 2.36 ;
        RECT  2.21 0.65 2.49 1.23 ;
        RECT  2.21 1.07 2.88 1.23 ;
        RECT  2.72 1.52 3.68 1.68 ;
        RECT  3.40 1.46 3.68 1.74 ;
        RECT  2.72 1.07 2.88 2.48 ;
        RECT  2.66 1.90 2.94 2.48 ;
        RECT  5.22 0.95 5.50 1.23 ;
        RECT  5.30 0.95 5.46 2.13 ;
        RECT  4.78 1.97 5.46 2.13 ;
        RECT  4.78 1.97 5.06 2.25 ;
        RECT  4.84 1.97 5.00 2.76 ;
        RECT  4.64 2.48 5.00 2.76 ;
    END
END NOR5SP4V1_0

MACRO NOR5SP2V1_0
    CLASS CORE ;
    FOREIGN NOR5SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 9.80  LAYER ME1  ;
        ANTENNADIFFAREA 4.79  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.34  LAYER ME1  ;
        ANTENNAMAXAREACAR 29.16  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.86 1.52 4.28 1.68 ;
        RECT  3.74 1.90 4.02 2.18 ;
        RECT  3.86 0.63 4.02 2.18 ;
        RECT  3.67 0.63 4.02 1.23 ;
        END
    END OUT
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.39 1.62 1.81 ;
        END
    END IN3
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.46 1.39 4.74 1.81 ;
        END
    END IN4
    PIN IN5
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.22 1.39 5.50 1.81 ;
        END
    END IN5
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 5.60 3.48 ;
        RECT  5.22 1.97 5.50 2.25 ;
        RECT  5.14 2.88 5.44 3.48 ;
        RECT  5.28 1.97 5.44 3.48 ;
        RECT  3.22 1.90 3.50 2.50 ;
        RECT  3.28 1.90 3.44 3.48 ;
        RECT  2.14 1.90 2.42 2.30 ;
        RECT  2.20 1.90 2.36 3.48 ;
        RECT  0.24 2.08 0.52 2.36 ;
        RECT  0.30 2.08 0.46 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 5.60 0.28 ;
        RECT  5.22 0.95 5.50 1.23 ;
        RECT  5.28 -0.28 5.44 1.23 ;
        RECT  5.14 -0.28 5.44 0.32 ;
        RECT  4.18 0.95 4.46 1.23 ;
        RECT  4.24 -0.28 4.40 1.23 ;
        RECT  3.15 0.63 3.43 1.23 ;
        RECT  3.21 -0.28 3.37 1.23 ;
        RECT  1.14 0.63 1.42 0.91 ;
        RECT  1.20 -0.28 1.36 0.91 ;
        RECT  0.10 0.63 0.38 0.91 ;
        RECT  0.16 -0.28 0.32 0.91 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.63 0.90 0.91 ;
        RECT  1.66 0.63 1.94 0.91 ;
        RECT  0.74 0.63 0.90 1.23 ;
        RECT  0.74 1.07 1.94 1.23 ;
        RECT  1.78 1.52 2.56 1.68 ;
        RECT  2.28 1.46 2.56 1.74 ;
        RECT  1.78 0.63 1.94 2.36 ;
        RECT  1.52 2.08 1.94 2.36 ;
        RECT  2.21 0.83 2.49 1.23 ;
        RECT  2.21 1.07 2.88 1.23 ;
        RECT  2.72 1.52 3.68 1.68 ;
        RECT  3.40 1.46 3.68 1.74 ;
        RECT  2.72 1.07 2.88 2.30 ;
        RECT  2.66 1.90 2.94 2.30 ;
        RECT  4.70 0.95 5.06 1.23 ;
        RECT  4.90 0.95 5.06 2.13 ;
        RECT  4.32 1.97 5.06 2.13 ;
        RECT  4.32 1.97 4.60 2.25 ;
        RECT  4.32 1.97 4.48 2.76 ;
        RECT  4.12 2.48 4.48 2.76 ;
    END
END NOR5SP2V1_0

MACRO NOR5SP1V1_0
    CLASS CORE ;
    FOREIGN NOR5SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN5
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.22 1.39 5.50 1.81 ;
        END
    END IN5
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.46 1.39 4.74 1.81 ;
        END
    END IN4
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 9.63  LAYER ME1  ;
        ANTENNADIFFAREA 4.14  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        ANTENNAMAXAREACAR 47.76  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.82 1.52 4.28 1.68 ;
        RECT  3.70 1.90 3.98 2.18 ;
        RECT  3.82 0.95 3.98 2.18 ;
        RECT  3.63 0.95 3.98 1.23 ;
        END
    END OUT
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.39 1.62 1.81 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 5.60 0.28 ;
        RECT  5.22 0.95 5.50 1.23 ;
        RECT  5.28 -0.28 5.44 1.23 ;
        RECT  5.14 -0.28 5.44 0.32 ;
        RECT  4.18 0.95 4.46 1.23 ;
        RECT  4.24 -0.28 4.40 1.23 ;
        RECT  3.11 0.95 3.39 1.23 ;
        RECT  3.17 -0.28 3.33 1.23 ;
        RECT  1.14 0.63 1.42 0.91 ;
        RECT  1.20 -0.28 1.36 0.91 ;
        RECT  0.10 0.63 0.38 0.91 ;
        RECT  0.16 -0.28 0.32 0.91 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 5.60 3.48 ;
        RECT  5.22 1.97 5.50 2.25 ;
        RECT  5.14 2.88 5.44 3.48 ;
        RECT  5.28 1.97 5.44 3.48 ;
        RECT  3.18 1.90 3.46 2.18 ;
        RECT  3.24 1.90 3.40 3.48 ;
        RECT  2.14 1.90 2.42 2.18 ;
        RECT  2.20 1.90 2.36 3.48 ;
        RECT  0.24 2.08 0.52 2.36 ;
        RECT  0.30 2.08 0.46 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.63 0.90 0.91 ;
        RECT  1.66 0.63 1.94 0.91 ;
        RECT  0.74 0.63 0.90 1.23 ;
        RECT  0.74 1.07 1.94 1.23 ;
        RECT  1.78 1.52 2.56 1.68 ;
        RECT  2.28 1.46 2.56 1.74 ;
        RECT  1.78 0.63 1.94 2.36 ;
        RECT  1.52 2.08 1.94 2.36 ;
        RECT  2.21 0.95 2.49 1.23 ;
        RECT  2.21 1.07 2.88 1.23 ;
        RECT  2.72 1.52 3.61 1.68 ;
        RECT  3.33 1.46 3.61 1.74 ;
        RECT  2.72 1.07 2.88 2.18 ;
        RECT  2.66 1.90 2.94 2.18 ;
        RECT  4.70 0.95 5.06 1.23 ;
        RECT  4.90 0.95 5.06 2.13 ;
        RECT  4.32 1.97 5.06 2.13 ;
        RECT  4.32 1.97 4.60 2.25 ;
        RECT  4.32 1.97 4.48 2.76 ;
        RECT  4.12 2.48 4.48 2.76 ;
    END
END NOR5SP1V1_0

MACRO NOR4SP8V1_0
    CLASS CORE ;
    FOREIGN NOR4SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.06 1.39 6.34 1.81 ;
        END
    END IN4
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.26 1.39 5.54 1.81 ;
        END
    END IN3
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 13.21  LAYER ME1  ;
        ANTENNADIFFAREA 7.30  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.91  LAYER ME1  ;
        ANTENNAMAXAREACAR 14.48  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.26 1.90 4.54 2.50 ;
        RECT  4.19 0.63 4.47 1.23 ;
        RECT  4.26 0.63 4.42 2.50 ;
        RECT  3.32 1.52 4.42 1.68 ;
        RECT  3.22 1.90 3.50 2.50 ;
        RECT  3.32 0.63 3.48 2.50 ;
        RECT  3.15 0.63 3.48 1.23 ;
        END
    END OUT
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 6.80 0.28 ;
        RECT  6.32 -0.28 6.62 0.32 ;
        RECT  6.26 0.95 6.54 1.23 ;
        RECT  6.32 -0.28 6.48 1.23 ;
        RECT  5.22 0.95 5.50 1.23 ;
        RECT  5.28 -0.28 5.44 1.23 ;
        RECT  4.71 0.63 4.99 1.23 ;
        RECT  4.77 -0.28 4.93 1.23 ;
        RECT  3.67 0.63 3.95 1.23 ;
        RECT  3.73 -0.28 3.89 1.23 ;
        RECT  2.59 0.53 2.87 1.23 ;
        RECT  2.65 -0.28 2.81 1.23 ;
        RECT  1.14 0.95 1.42 1.23 ;
        RECT  1.20 -0.28 1.36 1.23 ;
        RECT  0.10 0.95 0.38 1.23 ;
        RECT  0.16 -0.28 0.32 1.23 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 6.80 3.48 ;
        RECT  6.26 2.88 6.62 3.48 ;
        RECT  6.20 1.97 6.48 2.25 ;
        RECT  6.26 1.97 6.42 3.48 ;
        RECT  4.78 1.90 5.06 2.35 ;
        RECT  4.84 1.90 5.00 3.48 ;
        RECT  3.74 1.90 4.02 2.50 ;
        RECT  3.80 1.90 3.96 3.48 ;
        RECT  2.66 1.90 2.94 2.60 ;
        RECT  2.72 1.90 2.88 3.48 ;
        RECT  1.62 1.90 1.90 2.60 ;
        RECT  1.68 1.90 1.84 3.48 ;
        RECT  0.10 1.97 0.38 2.25 ;
        RECT  0.16 1.97 0.32 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.54 0.95 0.90 1.23 ;
        RECT  1.30 1.52 2.04 1.68 ;
        RECT  1.76 1.46 2.04 1.74 ;
        RECT  0.54 0.95 0.70 2.13 ;
        RECT  1.30 1.52 1.46 2.13 ;
        RECT  0.54 1.97 1.46 2.13 ;
        RECT  1.00 1.97 1.28 2.25 ;
        RECT  1.69 0.53 1.97 1.23 ;
        RECT  1.69 1.07 2.36 1.23 ;
        RECT  2.20 1.52 3.16 1.68 ;
        RECT  2.88 1.46 3.16 1.74 ;
        RECT  2.20 1.07 2.36 2.60 ;
        RECT  2.14 1.90 2.42 2.60 ;
        RECT  5.70 0.95 6.02 1.23 ;
        RECT  5.70 0.95 5.86 2.13 ;
        RECT  5.30 1.97 5.86 2.13 ;
        RECT  5.30 1.97 5.58 2.25 ;
        RECT  5.36 1.97 5.52 2.76 ;
        RECT  5.16 2.48 5.52 2.76 ;
    END
END NOR4SP8V1_0

MACRO NOR4SP4V1_0
    CLASS CORE ;
    FOREIGN NOR4SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.22 1.39 5.50 1.81 ;
        END
    END IN4
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.06 1.39 4.34 1.81 ;
        END
    END IN3
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 10.69  LAYER ME1  ;
        ANTENNADIFFAREA 5.25  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER ME1  ;
        ANTENNAMAXAREACAR 18.88  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.22 1.90 3.50 2.50 ;
        RECT  3.32 0.63 3.48 2.50 ;
        RECT  3.15 0.63 3.48 1.23 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 5.60 3.48 ;
        RECT  5.16 1.97 5.44 2.25 ;
        RECT  5.14 2.88 5.42 3.48 ;
        RECT  5.21 1.97 5.37 3.48 ;
        RECT  3.74 1.97 4.02 2.25 ;
        RECT  3.80 1.97 3.96 3.48 ;
        RECT  2.70 1.90 2.98 2.50 ;
        RECT  2.76 1.90 2.92 3.48 ;
        RECT  1.62 1.90 1.90 2.48 ;
        RECT  1.68 1.90 1.84 3.48 ;
        RECT  0.10 1.97 0.38 2.25 ;
        RECT  0.16 1.97 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 5.60 0.28 ;
        RECT  5.22 0.95 5.50 1.23 ;
        RECT  5.28 -0.28 5.44 1.23 ;
        RECT  5.14 -0.28 5.44 0.32 ;
        RECT  4.18 0.95 4.46 1.23 ;
        RECT  4.24 -0.28 4.40 1.23 ;
        RECT  3.67 0.63 3.95 1.23 ;
        RECT  3.73 -0.28 3.89 1.23 ;
        RECT  2.63 0.63 2.91 1.23 ;
        RECT  2.69 -0.28 2.85 1.23 ;
        RECT  1.14 0.95 1.42 1.23 ;
        RECT  1.20 -0.28 1.36 1.23 ;
        RECT  0.10 0.95 0.38 1.23 ;
        RECT  0.16 -0.28 0.32 1.23 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.54 0.95 0.90 1.23 ;
        RECT  1.30 1.52 2.04 1.68 ;
        RECT  1.76 1.46 2.04 1.74 ;
        RECT  0.54 0.95 0.70 2.13 ;
        RECT  1.30 1.52 1.46 2.13 ;
        RECT  0.54 1.97 1.46 2.13 ;
        RECT  1.00 1.97 1.28 2.25 ;
        RECT  1.69 0.65 1.97 1.23 ;
        RECT  1.69 1.07 2.36 1.23 ;
        RECT  2.20 1.52 3.16 1.68 ;
        RECT  2.88 1.46 3.16 1.74 ;
        RECT  2.20 1.07 2.36 2.48 ;
        RECT  2.14 1.90 2.42 2.48 ;
        RECT  4.66 0.95 4.98 1.23 ;
        RECT  4.66 0.95 4.82 2.13 ;
        RECT  4.26 1.97 4.82 2.13 ;
        RECT  4.26 1.97 4.54 2.25 ;
        RECT  4.32 1.97 4.48 2.76 ;
        RECT  4.12 2.48 4.48 2.76 ;
    END
END NOR4SP4V1_0

MACRO NOR4SP2V1_0
    CLASS CORE ;
    FOREIGN NOR4SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 9.24  LAYER ME1  ;
        ANTENNADIFFAREA 4.36  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.34  LAYER ME1  ;
        ANTENNAMAXAREACAR 27.51  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.22 1.90 3.50 2.18 ;
        RECT  3.32 0.63 3.48 2.18 ;
        RECT  3.15 0.63 3.48 1.23 ;
        END
    END OUT
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.46 1.39 4.74 1.81 ;
        END
    END IN4
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.66 1.39 3.94 1.81 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 5.20 0.28 ;
        RECT  4.74 -0.28 5.02 0.32 ;
        RECT  4.71 0.95 4.99 1.23 ;
        RECT  4.76 -0.28 4.92 1.23 ;
        RECT  3.67 0.95 3.95 1.23 ;
        RECT  3.72 -0.28 3.88 1.23 ;
        RECT  2.63 0.63 2.91 1.23 ;
        RECT  2.69 -0.28 2.85 1.23 ;
        RECT  1.14 0.95 1.42 1.23 ;
        RECT  1.20 -0.28 1.36 1.23 ;
        RECT  0.10 0.95 0.38 1.23 ;
        RECT  0.16 -0.28 0.32 1.23 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 5.20 3.48 ;
        RECT  4.69 2.88 5.02 3.48 ;
        RECT  4.64 1.97 4.92 2.25 ;
        RECT  4.69 1.97 4.85 3.48 ;
        RECT  2.70 1.90 2.98 2.50 ;
        RECT  2.76 1.90 2.92 3.48 ;
        RECT  1.62 1.90 1.90 2.30 ;
        RECT  1.68 1.90 1.84 3.48 ;
        RECT  0.10 1.97 0.38 2.25 ;
        RECT  0.16 1.97 0.32 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.54 0.95 0.90 1.23 ;
        RECT  1.30 1.52 2.04 1.68 ;
        RECT  1.76 1.46 2.04 1.74 ;
        RECT  0.54 0.95 0.70 2.13 ;
        RECT  1.30 1.52 1.46 2.13 ;
        RECT  0.54 1.97 1.46 2.13 ;
        RECT  1.00 1.97 1.28 2.25 ;
        RECT  1.69 0.83 1.97 1.23 ;
        RECT  1.69 1.07 2.36 1.23 ;
        RECT  2.20 1.52 3.16 1.68 ;
        RECT  2.88 1.46 3.16 1.74 ;
        RECT  2.20 1.07 2.36 2.30 ;
        RECT  2.14 1.90 2.42 2.30 ;
        RECT  4.14 0.95 4.47 1.23 ;
        RECT  4.14 0.95 4.30 2.13 ;
        RECT  3.74 1.97 4.30 2.13 ;
        RECT  3.74 1.97 4.02 2.25 ;
        RECT  3.80 1.97 3.96 2.76 ;
        RECT  3.60 2.48 3.96 2.76 ;
    END
END NOR4SP2V1_0

MACRO NOR4SP1V1_0
    CLASS CORE ;
    FOREIGN NOR4SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.66 1.39 3.94 1.81 ;
        END
    END IN3
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.46 1.39 4.74 1.81 ;
        END
    END IN4
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 9.03  LAYER ME1  ;
        ANTENNADIFFAREA 3.72  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        ANTENNAMAXAREACAR 44.80  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.18 1.97 3.48 2.25 ;
        RECT  3.32 0.95 3.48 2.25 ;
        RECT  3.11 0.95 3.48 1.23 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 5.20 3.48 ;
        RECT  4.67 2.88 5.02 3.48 ;
        RECT  4.61 1.97 4.89 2.25 ;
        RECT  4.67 1.97 4.83 3.48 ;
        RECT  2.66 1.97 2.94 2.25 ;
        RECT  2.72 1.97 2.88 3.48 ;
        RECT  1.62 1.97 1.90 2.25 ;
        RECT  1.68 1.97 1.84 3.48 ;
        RECT  0.10 1.97 0.38 2.25 ;
        RECT  0.16 1.97 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 5.20 0.28 ;
        RECT  4.74 -0.28 5.02 0.32 ;
        RECT  4.68 0.95 4.96 1.23 ;
        RECT  4.74 -0.28 4.90 1.23 ;
        RECT  3.64 0.95 3.92 1.23 ;
        RECT  3.70 -0.28 3.86 1.23 ;
        RECT  2.59 0.95 2.87 1.23 ;
        RECT  2.65 -0.28 2.81 1.23 ;
        RECT  1.14 0.95 1.42 1.23 ;
        RECT  1.20 -0.28 1.36 1.23 ;
        RECT  0.10 0.95 0.38 1.23 ;
        RECT  0.16 -0.28 0.32 1.23 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.54 0.95 0.90 1.23 ;
        RECT  1.30 1.52 2.04 1.68 ;
        RECT  1.76 1.46 2.04 1.74 ;
        RECT  0.54 0.95 0.70 2.13 ;
        RECT  1.30 1.52 1.46 2.13 ;
        RECT  0.54 1.97 1.46 2.13 ;
        RECT  1.00 1.97 1.28 2.25 ;
        RECT  1.69 0.95 1.97 1.23 ;
        RECT  1.69 1.07 2.36 1.23 ;
        RECT  2.20 1.52 3.08 1.68 ;
        RECT  2.80 1.46 3.08 1.74 ;
        RECT  2.20 1.07 2.36 2.25 ;
        RECT  2.14 1.97 2.42 2.25 ;
        RECT  4.14 0.95 4.44 1.23 ;
        RECT  4.14 0.95 4.30 2.13 ;
        RECT  3.71 1.97 4.30 2.13 ;
        RECT  3.71 1.97 3.99 2.25 ;
        RECT  3.71 1.97 3.87 2.69 ;
        RECT  3.57 2.41 3.87 2.69 ;
    END
END NOR4SP1V1_0

MACRO NOR3SP8V1_0
    CLASS CORE ;
    FOREIGN NOR3SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.58  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.46 1.39 2.74 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.58  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN1
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.58  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.86 1.39 5.14 1.81 ;
        END
    END IN3
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 12.89  LAYER ME1  ;
        ANTENNADIFFAREA 8.87  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.30 1.97 6.58 2.25 ;
        RECT  0.74 1.07 6.58 1.23 ;
        RECT  6.30 0.95 6.58 1.23 ;
        RECT  5.26 1.97 6.58 2.13 ;
        RECT  5.26 1.97 5.54 2.25 ;
        RECT  5.26 0.95 5.54 1.23 ;
        RECT  5.32 0.95 5.48 2.25 ;
        RECT  3.74 0.79 4.02 1.23 ;
        RECT  2.70 0.79 2.98 1.23 ;
        RECT  1.66 0.79 1.94 1.23 ;
        RECT  0.62 0.79 0.90 1.07 ;
        END
    END OUT
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 7.20 0.28 ;
        RECT  6.82 0.63 7.10 0.91 ;
        RECT  6.88 -0.28 7.04 0.91 ;
        RECT  6.74 -0.28 7.04 0.32 ;
        RECT  5.78 0.63 6.06 0.91 ;
        RECT  5.84 -0.28 6.00 0.91 ;
        RECT  4.74 0.63 5.02 0.91 ;
        RECT  4.80 -0.28 4.96 0.91 ;
        RECT  4.26 0.63 4.54 0.91 ;
        RECT  4.32 -0.28 4.48 0.91 ;
        RECT  3.22 0.63 3.50 0.91 ;
        RECT  3.28 -0.28 3.44 0.91 ;
        RECT  2.18 0.63 2.46 0.91 ;
        RECT  2.24 -0.28 2.40 0.91 ;
        RECT  1.14 0.63 1.42 0.91 ;
        RECT  1.20 -0.28 1.36 0.91 ;
        RECT  0.10 0.63 0.38 0.91 ;
        RECT  0.16 -0.28 0.32 0.91 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 7.20 3.48 ;
        RECT  6.74 2.88 7.02 3.48 ;
        RECT  1.66 2.29 1.94 2.57 ;
        RECT  1.72 2.29 1.88 3.48 ;
        RECT  0.62 2.29 0.90 2.57 ;
        RECT  0.68 2.29 0.84 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.10 1.97 4.54 2.13 ;
        RECT  0.10 1.97 0.38 2.25 ;
        RECT  1.14 1.97 1.42 2.25 ;
        RECT  2.18 1.97 2.46 2.25 ;
        RECT  3.22 1.97 3.50 2.25 ;
        RECT  4.26 1.97 4.54 2.25 ;
        RECT  2.70 2.29 2.98 2.57 ;
        RECT  3.74 2.29 4.02 2.57 ;
        RECT  4.74 2.29 5.02 2.57 ;
        RECT  5.78 2.29 6.06 2.57 ;
        RECT  6.82 2.29 7.10 2.57 ;
        RECT  2.70 2.41 7.10 2.57 ;
    END
END NOR3SP8V1_0

MACRO NOR3SP4V1_0
    CLASS CORE ;
    FOREIGN NOR3SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.29  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.06 1.39 2.34 1.81 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.29  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.66 1.39 3.94 1.81 ;
        END
    END IN3
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.29  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN1
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 7.48  LAYER ME1  ;
        ANTENNADIFFAREA 5.09  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.18 2.05 3.48 2.33 ;
        RECT  3.32 0.86 3.48 2.33 ;
        RECT  0.74 0.98 3.48 1.14 ;
        RECT  3.18 0.86 3.48 1.14 ;
        RECT  1.66 0.70 1.94 1.14 ;
        RECT  0.62 0.70 0.90 0.98 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.40 3.48 ;
        RECT  3.94 2.88 4.22 3.48 ;
        RECT  0.62 2.37 0.90 2.65 ;
        RECT  0.68 2.37 0.84 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.40 0.28 ;
        RECT  3.76 -0.28 4.22 0.32 ;
        RECT  3.70 0.54 3.98 0.82 ;
        RECT  3.76 -0.28 3.92 0.82 ;
        RECT  2.66 0.54 2.94 0.82 ;
        RECT  2.72 -0.28 2.88 0.82 ;
        RECT  2.18 0.54 2.46 0.82 ;
        RECT  2.24 -0.28 2.40 0.82 ;
        RECT  1.14 0.54 1.42 0.82 ;
        RECT  1.20 -0.28 1.36 0.82 ;
        RECT  0.10 0.54 0.38 0.82 ;
        RECT  0.16 -0.28 0.32 0.82 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.10 2.05 2.46 2.21 ;
        RECT  0.10 2.05 0.38 2.33 ;
        RECT  1.14 2.05 1.42 2.33 ;
        RECT  2.18 2.05 2.46 2.33 ;
        RECT  1.66 2.37 1.94 2.65 ;
        RECT  2.66 2.37 2.94 2.65 ;
        RECT  3.70 2.37 3.98 2.65 ;
        RECT  1.66 2.49 3.98 2.65 ;
    END
END NOR3SP4V1_0

MACRO NOR3SP2V1_0
    CLASS CORE ;
    FOREIGN NOR3SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 2.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 3.16  LAYER ME1  ;
        ANTENNADIFFAREA 2.51  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.52 2.05 2.28 2.21 ;
        RECT  2.12 0.98 2.28 2.21 ;
        RECT  0.74 0.98 2.28 1.14 ;
        RECT  1.66 0.70 1.94 1.14 ;
        RECT  1.52 2.05 1.80 2.65 ;
        RECT  0.62 0.70 0.90 0.98 ;
        END
    END OUT
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.14  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.14  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.28 1.39 1.58 1.81 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.14  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.82 1.39 1.12 1.81 ;
        END
    END IN2
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 2.40 0.28 ;
        RECT  1.94 -0.28 2.22 0.32 ;
        RECT  1.14 0.54 1.42 0.82 ;
        RECT  1.20 -0.28 1.36 0.82 ;
        RECT  0.10 0.54 0.38 0.82 ;
        RECT  0.16 -0.28 0.32 0.82 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 2.40 3.48 ;
        RECT  1.94 2.88 2.22 3.48 ;
        RECT  0.24 2.05 0.52 2.65 ;
        RECT  0.30 2.05 0.46 3.48 ;
        END
    END VDD!
END NOR3SP2V1_0

MACRO NOR3SP1V1_0
    CLASS CORE ;
    FOREIGN NOR3SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 2.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.10  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.10  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.82 1.44 1.10 1.86 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.10  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.44 1.58 1.86 ;
        END
    END IN3
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 3.18  LAYER ME1  ;
        ANTENNADIFFAREA 1.99  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.78 1.12 1.94 2.28 ;
        RECT  1.66 0.64 1.94 0.92 ;
        RECT  1.66 0.64 1.82 1.28 ;
        RECT  1.52 2.12 1.80 2.68 ;
        RECT  0.74 1.12 1.94 1.28 ;
        RECT  0.74 0.64 0.90 1.28 ;
        RECT  0.62 0.64 0.90 0.92 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 2.40 3.48 ;
        RECT  1.94 2.88 2.22 3.48 ;
        RECT  0.24 2.12 0.52 2.68 ;
        RECT  0.30 2.12 0.46 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 2.40 0.28 ;
        RECT  1.94 -0.28 2.22 0.32 ;
        RECT  1.14 0.64 1.42 0.92 ;
        RECT  1.20 -0.28 1.36 0.92 ;
        RECT  0.10 0.64 0.38 0.92 ;
        RECT  0.16 -0.28 0.32 0.92 ;
        END
    END GND!
END NOR3SP1V1_0

MACRO NOR2SP8V1_0
    CLASS CORE ;
    FOREIGN NOR2SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.59  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.59  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.39 1.46 2.81 1.74 ;
        END
    END IN2
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 8.39  LAYER ME1  ;
        ANTENNADIFFAREA 5.92  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.66 1.08 4.06 1.24 ;
        RECT  3.78 0.96 4.06 1.24 ;
        RECT  2.74 0.96 3.02 1.24 ;
        RECT  1.70 1.90 1.98 2.18 ;
        RECT  1.70 0.96 1.98 1.24 ;
        RECT  0.66 1.92 1.98 2.08 ;
        RECT  0.86 1.46 1.14 1.74 ;
        RECT  0.92 1.08 1.08 2.08 ;
        RECT  0.66 1.92 0.94 2.20 ;
        RECT  0.66 0.96 0.94 1.24 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.80 3.48 ;
        RECT  4.34 2.88 4.62 3.48 ;
        RECT  3.78 2.24 4.06 2.52 ;
        RECT  3.84 2.24 4.00 3.48 ;
        RECT  2.74 2.24 3.02 2.52 ;
        RECT  2.80 2.24 2.96 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.80 0.28 ;
        RECT  4.34 -0.28 4.62 0.32 ;
        RECT  4.30 0.64 4.58 0.92 ;
        RECT  4.36 -0.28 4.52 0.92 ;
        RECT  3.26 0.64 3.54 0.92 ;
        RECT  3.32 -0.28 3.48 0.92 ;
        RECT  2.22 0.64 2.50 0.92 ;
        RECT  2.28 -0.28 2.44 0.92 ;
        RECT  1.18 0.64 1.46 0.92 ;
        RECT  1.24 -0.28 1.40 0.92 ;
        RECT  0.14 0.64 0.42 0.92 ;
        RECT  0.20 -0.28 0.36 0.92 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  2.34 1.90 4.58 2.06 ;
        RECT  3.26 1.90 3.54 2.18 ;
        RECT  4.30 1.90 4.58 2.18 ;
        RECT  0.14 2.24 0.42 2.52 ;
        RECT  1.18 2.24 1.46 2.52 ;
        RECT  2.22 2.24 2.50 2.52 ;
        RECT  2.34 1.90 2.50 2.52 ;
        RECT  0.14 2.36 2.50 2.52 ;
    END
END NOR2SP8V1_0

MACRO NOR2SP4V1_0
    CLASS CORE ;
    FOREIGN NOR2SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 2.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 4.23  LAYER ME1  ;
        ANTENNADIFFAREA 3.56  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.66 1.08 1.98 1.24 ;
        RECT  1.70 0.96 1.98 1.24 ;
        RECT  0.92 1.08 1.08 2.11 ;
        RECT  0.66 1.90 0.94 2.18 ;
        RECT  0.66 0.96 0.94 1.24 ;
        END
    END OUT
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.29  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.29  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.99 1.46 2.41 1.74 ;
        END
    END IN2
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 2.80 3.48 ;
        RECT  2.34 2.88 2.62 3.48 ;
        RECT  1.70 2.24 1.98 2.52 ;
        RECT  1.76 2.24 1.92 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 2.80 0.28 ;
        RECT  2.28 -0.28 2.62 0.32 ;
        RECT  2.22 0.64 2.50 0.92 ;
        RECT  2.28 -0.28 2.44 0.92 ;
        RECT  1.18 0.64 1.46 0.92 ;
        RECT  1.24 -0.28 1.40 0.92 ;
        RECT  0.14 0.64 0.42 0.92 ;
        RECT  0.20 -0.28 0.36 0.92 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  1.30 1.92 2.50 2.08 ;
        RECT  2.22 1.90 2.50 2.18 ;
        RECT  0.14 2.24 0.42 2.52 ;
        RECT  1.18 2.24 1.46 2.52 ;
        RECT  1.30 1.92 1.46 2.52 ;
        RECT  0.14 2.36 1.46 2.52 ;
    END
END NOR2SP4V1_0

MACRO NOR2SP2V1_0
    CLASS CORE ;
    FOREIGN NOR2SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 1.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.14  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.42 1.44 0.70 1.86 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.14  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.90 1.44 1.18 1.86 ;
        END
    END IN2
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 2.29  LAYER ME1  ;
        ANTENNADIFFAREA 1.86  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.34 1.12 1.50 2.18 ;
        RECT  1.11 2.02 1.39 2.62 ;
        RECT  0.64 1.12 1.50 1.28 ;
        RECT  0.64 0.95 0.92 1.28 ;
        END
    END OUT
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 1.60 0.28 ;
        RECT  1.16 0.63 1.44 0.91 ;
        RECT  1.14 -0.28 1.42 0.32 ;
        RECT  1.22 -0.28 1.38 0.91 ;
        RECT  0.12 0.63 0.40 0.91 ;
        RECT  0.18 -0.28 0.34 0.91 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 1.60 3.48 ;
        RECT  1.14 2.88 1.42 3.48 ;
        RECT  0.21 2.02 0.49 2.62 ;
        RECT  0.27 2.02 0.43 3.48 ;
        END
    END VDD!
END NOR2SP2V1_0

MACRO NOR2SP1V1_0
    CLASS CORE ;
    FOREIGN NOR2SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 1.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.42 1.44 0.70 1.86 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.90 1.44 1.18 1.86 ;
        END
    END IN2
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 2.25  LAYER ME1  ;
        ANTENNADIFFAREA 1.21  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.11 2.02 1.50 2.30 ;
        RECT  1.34 1.12 1.50 2.30 ;
        RECT  0.76 1.12 1.50 1.28 ;
        RECT  0.76 0.63 0.92 1.28 ;
        RECT  0.64 0.63 0.92 0.91 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 1.60 3.48 ;
        RECT  1.14 2.88 1.42 3.48 ;
        RECT  0.21 2.02 0.49 2.30 ;
        RECT  0.27 2.02 0.43 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 1.60 0.28 ;
        RECT  1.16 0.63 1.44 0.91 ;
        RECT  1.14 -0.28 1.42 0.32 ;
        RECT  1.22 -0.28 1.38 0.91 ;
        RECT  0.12 0.63 0.40 0.91 ;
        RECT  0.18 -0.28 0.34 0.91 ;
        END
    END GND!
END NOR2SP1V1_0

MACRO NOR2SP16V1_0
    CLASS CORE ;
    FOREIGN NOR2SP16V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.17  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.17  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.39 1.46 4.81 1.74 ;
        END
    END IN2
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 16.12  LAYER ME1  ;
        ANTENNADIFFAREA 11.23  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.66 1.08 8.22 1.24 ;
        RECT  7.94 0.96 8.22 1.24 ;
        RECT  6.90 0.96 7.18 1.24 ;
        RECT  5.86 0.96 6.14 1.24 ;
        RECT  4.82 0.96 5.10 1.24 ;
        RECT  3.78 1.90 4.06 2.18 ;
        RECT  3.78 0.96 4.06 1.24 ;
        RECT  0.66 1.92 4.06 2.08 ;
        RECT  2.74 1.90 3.02 2.18 ;
        RECT  2.74 0.96 3.02 1.24 ;
        RECT  1.70 1.90 1.98 2.18 ;
        RECT  1.70 0.96 1.98 1.24 ;
        RECT  0.92 1.08 1.08 2.08 ;
        RECT  0.66 1.92 0.94 2.20 ;
        RECT  0.66 0.96 0.94 1.24 ;
        END
    END OUT
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 9.20 0.28 ;
        RECT  8.52 -0.28 9.02 0.32 ;
        RECT  8.46 0.64 8.74 0.92 ;
        RECT  8.52 -0.28 8.68 0.92 ;
        RECT  7.42 0.64 7.70 0.92 ;
        RECT  7.48 -0.28 7.64 0.92 ;
        RECT  6.38 0.64 6.66 0.92 ;
        RECT  6.44 -0.28 6.60 0.92 ;
        RECT  5.34 0.64 5.62 0.92 ;
        RECT  5.40 -0.28 5.56 0.92 ;
        RECT  4.30 0.64 4.58 0.92 ;
        RECT  4.36 -0.28 4.52 0.92 ;
        RECT  3.26 0.64 3.54 0.92 ;
        RECT  3.32 -0.28 3.48 0.92 ;
        RECT  2.22 0.64 2.50 0.92 ;
        RECT  2.28 -0.28 2.44 0.92 ;
        RECT  1.18 0.64 1.46 0.92 ;
        RECT  1.24 -0.28 1.40 0.92 ;
        RECT  0.14 0.64 0.42 0.92 ;
        RECT  0.20 -0.28 0.36 0.92 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 9.20 3.48 ;
        RECT  8.74 2.88 9.02 3.48 ;
        RECT  7.94 2.24 8.22 2.52 ;
        RECT  8.00 2.24 8.16 3.48 ;
        RECT  6.90 2.24 7.18 2.52 ;
        RECT  6.96 2.24 7.12 3.48 ;
        RECT  5.86 2.24 6.14 2.52 ;
        RECT  5.92 2.24 6.08 3.48 ;
        RECT  4.82 2.24 5.10 2.52 ;
        RECT  4.88 2.24 5.04 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  4.42 1.92 8.74 2.08 ;
        RECT  5.34 1.90 5.62 2.18 ;
        RECT  6.38 1.90 6.66 2.18 ;
        RECT  7.42 1.90 7.70 2.18 ;
        RECT  8.46 1.90 8.74 2.18 ;
        RECT  0.14 2.24 0.42 2.52 ;
        RECT  1.18 2.24 1.46 2.52 ;
        RECT  2.22 2.24 2.50 2.52 ;
        RECT  3.26 2.24 3.54 2.52 ;
        RECT  4.30 2.24 4.58 2.52 ;
        RECT  4.42 1.92 4.58 2.52 ;
        RECT  0.14 2.36 4.58 2.52 ;
    END
END NOR2SP16V1_0

MACRO NAND8SP8V1_0
    CLASS CORE ;
    FOREIGN NAND8SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN8
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.46 1.39 8.74 1.81 ;
        END
    END IN8
    PIN IN7
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.72 1.39 8.04 1.81 ;
        END
    END IN7
    PIN IN6
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.28 1.39 7.56 1.81 ;
        END
    END IN6
    PIN IN5
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.80 1.39 7.08 1.81 ;
        END
    END IN5
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.39 0.68 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.88 1.39 1.16 1.81 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.32 1.46 1.74 1.74 ;
        END
    END IN3
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.00 1.39 2.28 1.81 ;
        END
    END IN4
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 16.70  LAYER ME1  ;
        ANTENNADIFFAREA 8.95  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.89  LAYER ME1  ;
        ANTENNAMAXAREACAR 18.70  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.39 0.66 5.68 1.24 ;
        RECT  5.26 1.84 5.55 2.42 ;
        RECT  5.39 0.66 5.55 2.42 ;
        RECT  4.46 1.52 5.55 1.68 ;
        RECT  4.36 0.66 4.64 1.24 ;
        RECT  4.46 0.66 4.62 2.00 ;
        RECT  4.22 1.84 4.50 2.42 ;
        END
    END OUT
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 9.20 0.28 ;
        RECT  8.46 -0.28 9.02 0.32 ;
        RECT  8.40 0.63 8.68 0.91 ;
        RECT  8.46 -0.28 8.62 0.91 ;
        RECT  5.92 0.66 6.20 1.24 ;
        RECT  5.98 -0.28 6.14 1.24 ;
        RECT  4.88 0.66 5.16 1.24 ;
        RECT  4.94 -0.28 5.10 1.24 ;
        RECT  3.80 0.54 4.08 1.24 ;
        RECT  3.86 -0.28 4.02 1.24 ;
        RECT  2.76 0.54 3.04 1.24 ;
        RECT  2.82 -0.28 2.98 1.24 ;
        RECT  1.96 0.75 2.24 1.03 ;
        RECT  2.02 -0.28 2.18 1.03 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 9.20 3.48 ;
        RECT  8.66 2.88 9.02 3.48 ;
        RECT  8.60 2.29 8.88 2.57 ;
        RECT  8.66 2.29 8.82 3.48 ;
        RECT  7.56 2.29 7.84 2.57 ;
        RECT  7.62 2.29 7.78 3.48 ;
        RECT  6.52 2.29 6.80 2.57 ;
        RECT  6.58 2.29 6.74 3.48 ;
        RECT  5.78 1.84 6.06 2.42 ;
        RECT  5.84 1.84 6.00 3.48 ;
        RECT  4.74 2.14 5.02 2.42 ;
        RECT  4.80 2.14 4.96 3.48 ;
        RECT  3.66 1.84 3.94 2.54 ;
        RECT  3.72 1.84 3.88 3.48 ;
        RECT  1.66 2.29 1.94 2.57 ;
        RECT  1.72 2.29 1.88 3.48 ;
        RECT  0.62 2.29 0.90 2.57 ;
        RECT  0.68 2.29 0.84 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.08 0.75 0.58 1.03 ;
        RECT  2.44 1.40 2.88 1.68 ;
        RECT  0.08 0.75 0.24 2.13 ;
        RECT  2.44 1.40 2.60 2.13 ;
        RECT  0.08 1.97 2.60 2.13 ;
        RECT  0.16 1.97 0.32 2.57 ;
        RECT  1.20 1.97 1.36 2.57 ;
        RECT  2.24 1.97 2.40 2.57 ;
        RECT  0.10 2.29 0.38 2.57 ;
        RECT  1.14 2.29 1.42 2.57 ;
        RECT  2.18 2.29 2.46 2.57 ;
        RECT  3.20 0.54 3.56 1.24 ;
        RECT  3.20 1.46 4.30 1.62 ;
        RECT  4.02 1.40 4.30 1.68 ;
        RECT  3.20 0.54 3.36 2.00 ;
        RECT  2.76 1.84 3.36 2.00 ;
        RECT  2.76 1.84 3.04 2.54 ;
        RECT  6.74 0.63 7.02 0.91 ;
        RECT  6.36 0.75 7.02 0.91 ;
        RECT  6.20 1.46 6.52 1.74 ;
        RECT  6.36 0.75 6.52 2.13 ;
        RECT  6.36 1.97 8.36 2.13 ;
        RECT  7.16 1.97 7.32 2.57 ;
        RECT  7.04 2.29 7.32 2.57 ;
        RECT  8.20 1.97 8.36 2.57 ;
        RECT  8.08 2.29 8.36 2.57 ;
    END
END NAND8SP8V1_0

MACRO NAND8SP4V1_0
    CLASS CORE ;
    FOREIGN NAND8SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN8
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.28 1.39 7.56 1.81 ;
        END
    END IN8
    PIN IN7
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.80 1.39 7.08 1.81 ;
        END
    END IN7
    PIN IN6
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.10 1.39 6.38 1.81 ;
        END
    END IN6
    PIN IN5
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.62 1.39 5.90 1.81 ;
        END
    END IN5
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.39 0.68 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.88 1.39 1.16 1.81 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.32 1.46 1.74 1.74 ;
        END
    END IN3
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.00 1.39 2.28 1.81 ;
        END
    END IN4
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 13.76  LAYER ME1  ;
        ANTENNADIFFAREA 7.12  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.56  LAYER ME1  ;
        ANTENNAMAXAREACAR 24.72  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.46 1.52 4.68 1.68 ;
        RECT  4.46 0.66 4.62 2.00 ;
        RECT  4.18 1.84 4.46 2.42 ;
        RECT  4.32 0.66 4.62 1.24 ;
        END
    END OUT
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 8.00 0.28 ;
        RECT  7.38 -0.28 7.82 0.32 ;
        RECT  7.32 0.63 7.60 0.91 ;
        RECT  7.38 -0.28 7.54 0.91 ;
        RECT  4.84 0.66 5.12 1.24 ;
        RECT  4.90 -0.28 5.06 1.24 ;
        RECT  3.80 0.66 4.08 1.24 ;
        RECT  3.86 -0.28 4.02 1.24 ;
        RECT  2.76 0.66 3.04 1.24 ;
        RECT  2.82 -0.28 2.98 1.24 ;
        RECT  1.96 0.75 2.24 1.03 ;
        RECT  2.02 -0.28 2.18 1.03 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 8.00 3.48 ;
        RECT  7.54 2.88 7.82 3.48 ;
        RECT  7.52 2.29 7.80 2.57 ;
        RECT  7.58 2.29 7.74 3.48 ;
        RECT  6.48 2.29 6.76 2.57 ;
        RECT  6.54 2.29 6.70 3.48 ;
        RECT  5.44 2.29 5.72 2.57 ;
        RECT  5.50 2.29 5.66 3.48 ;
        RECT  4.70 2.14 4.98 2.42 ;
        RECT  4.76 2.14 4.92 3.48 ;
        RECT  3.66 1.84 3.94 2.42 ;
        RECT  3.72 1.84 3.88 3.48 ;
        RECT  1.66 2.29 1.94 2.57 ;
        RECT  1.72 2.29 1.88 3.48 ;
        RECT  0.62 2.29 0.90 2.57 ;
        RECT  0.68 2.29 0.84 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.08 0.75 0.58 1.03 ;
        RECT  2.44 1.40 2.88 1.68 ;
        RECT  0.08 0.75 0.24 2.13 ;
        RECT  2.44 1.40 2.60 2.13 ;
        RECT  0.08 1.97 2.60 2.13 ;
        RECT  0.16 1.97 0.32 2.57 ;
        RECT  1.20 1.97 1.36 2.57 ;
        RECT  2.24 1.97 2.40 2.57 ;
        RECT  0.10 2.29 0.38 2.57 ;
        RECT  1.14 2.29 1.42 2.57 ;
        RECT  2.18 2.29 2.46 2.57 ;
        RECT  3.20 0.66 3.56 1.24 ;
        RECT  3.20 1.46 4.28 1.62 ;
        RECT  4.00 1.40 4.28 1.68 ;
        RECT  3.20 0.66 3.36 2.00 ;
        RECT  2.76 1.84 3.36 2.00 ;
        RECT  2.76 1.84 3.04 2.42 ;
        RECT  5.66 0.63 5.94 0.91 ;
        RECT  5.28 0.75 5.94 0.91 ;
        RECT  5.12 1.46 5.44 1.74 ;
        RECT  5.28 0.75 5.44 2.13 ;
        RECT  5.28 1.97 7.28 2.13 ;
        RECT  6.08 1.97 6.24 2.57 ;
        RECT  5.96 2.29 6.24 2.57 ;
        RECT  7.12 1.97 7.28 2.57 ;
        RECT  7.00 2.29 7.28 2.57 ;
    END
END NAND8SP4V1_0

MACRO NAND8SP2V1_0
    CLASS CORE ;
    FOREIGN NAND8SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN8
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.92 1.39 7.22 1.81 ;
        END
    END IN8
    PIN IN7
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.46 1.39 6.74 1.81 ;
        END
    END IN7
    PIN IN6
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.72 1.39 6.04 1.81 ;
        END
    END IN6
    PIN IN5
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.26 1.39 5.54 1.81 ;
        END
    END IN5
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 12.87  LAYER ME1  ;
        ANTENNADIFFAREA 6.09  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.34  LAYER ME1  ;
        ANTENNAMAXAREACAR 38.31  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.46 1.52 4.68 1.68 ;
        RECT  4.36 0.64 4.64 1.24 ;
        RECT  4.46 0.64 4.62 2.00 ;
        RECT  4.22 1.84 4.50 2.44 ;
        END
    END OUT
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.00 1.39 2.28 1.81 ;
        END
    END IN4
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.32 1.46 1.74 1.74 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.88 1.39 1.16 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.39 0.68 1.81 ;
        END
    END IN1
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 7.60 0.28 ;
        RECT  7.04 -0.28 7.42 0.32 ;
        RECT  6.98 0.63 7.26 0.91 ;
        RECT  7.04 -0.28 7.20 0.91 ;
        RECT  3.84 0.64 4.12 1.24 ;
        RECT  3.90 -0.28 4.06 1.24 ;
        RECT  2.76 0.84 3.04 1.24 ;
        RECT  2.82 -0.28 2.98 1.24 ;
        RECT  1.96 0.75 2.24 1.03 ;
        RECT  2.02 -0.28 2.18 1.03 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 7.60 3.48 ;
        RECT  7.18 2.29 7.46 2.57 ;
        RECT  7.14 2.88 7.42 3.48 ;
        RECT  7.24 2.29 7.40 3.48 ;
        RECT  6.14 2.29 6.42 2.57 ;
        RECT  6.20 2.29 6.36 3.48 ;
        RECT  5.10 2.29 5.38 2.57 ;
        RECT  5.16 2.29 5.32 3.48 ;
        RECT  3.70 1.84 3.98 2.44 ;
        RECT  3.76 1.84 3.92 3.48 ;
        RECT  1.66 2.29 1.94 2.57 ;
        RECT  1.72 2.29 1.88 3.48 ;
        RECT  0.62 2.29 0.90 2.57 ;
        RECT  0.68 2.29 0.84 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.08 0.75 0.58 1.03 ;
        RECT  2.44 1.40 2.88 1.68 ;
        RECT  0.08 0.75 0.24 2.13 ;
        RECT  2.44 1.40 2.60 2.13 ;
        RECT  0.08 1.97 2.60 2.13 ;
        RECT  0.16 1.97 0.32 2.57 ;
        RECT  1.20 1.97 1.36 2.57 ;
        RECT  2.24 1.97 2.40 2.57 ;
        RECT  0.10 2.29 0.38 2.57 ;
        RECT  1.14 2.29 1.42 2.57 ;
        RECT  2.18 2.29 2.46 2.57 ;
        RECT  3.20 0.84 3.56 1.24 ;
        RECT  3.20 1.46 4.30 1.62 ;
        RECT  4.02 1.40 4.30 1.68 ;
        RECT  3.20 0.84 3.36 2.00 ;
        RECT  2.76 1.84 3.36 2.00 ;
        RECT  2.76 1.84 3.04 2.24 ;
        RECT  5.32 0.63 5.60 0.91 ;
        RECT  4.90 0.75 5.60 0.91 ;
        RECT  4.90 0.75 5.06 2.13 ;
        RECT  4.78 1.97 6.94 2.13 ;
        RECT  4.78 1.97 4.94 2.44 ;
        RECT  4.66 2.16 4.94 2.44 ;
        RECT  5.74 1.97 5.90 2.57 ;
        RECT  5.62 2.29 5.90 2.57 ;
        RECT  6.78 1.97 6.94 2.57 ;
        RECT  6.66 2.29 6.94 2.57 ;
    END
END NAND8SP2V1_0

MACRO NAND8SP1V1_0
    CLASS CORE ;
    FOREIGN NAND8SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN6
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.66 1.39 5.94 1.81 ;
        END
    END IN6
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.39 0.68 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.88 1.39 1.16 1.81 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.32 1.46 1.74 1.74 ;
        END
    END IN3
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.00 1.39 2.28 1.81 ;
        END
    END IN4
    PIN IN5
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.86 1.39 5.14 1.81 ;
        END
    END IN5
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 12.80  LAYER ME1  ;
        ANTENNADIFFAREA 5.34  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        ANTENNAMAXAREACAR 63.50  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.18 1.84 4.68 2.00 ;
        RECT  4.52 0.96 4.68 2.00 ;
        RECT  4.32 0.96 4.68 1.24 ;
        RECT  4.18 1.84 4.46 2.12 ;
        END
    END OUT
    PIN IN7
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.10 1.39 6.42 1.81 ;
        END
    END IN7
    PIN IN8
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.90 1.39 7.18 1.81 ;
        END
    END IN8
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 7.60 0.28 ;
        RECT  7.14 -0.28 7.42 0.32 ;
        RECT  6.70 0.63 6.98 0.91 ;
        RECT  6.76 -0.28 6.92 0.91 ;
        RECT  3.80 0.96 4.08 1.24 ;
        RECT  3.86 -0.28 4.02 1.24 ;
        RECT  2.76 0.96 3.04 1.24 ;
        RECT  2.82 -0.28 2.98 1.24 ;
        RECT  1.96 0.75 2.24 1.03 ;
        RECT  2.02 -0.28 2.18 1.03 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 7.60 3.48 ;
        RECT  6.96 2.88 7.42 3.48 ;
        RECT  6.90 2.29 7.18 2.57 ;
        RECT  6.96 2.29 7.12 3.48 ;
        RECT  5.86 2.29 6.14 2.57 ;
        RECT  5.92 2.29 6.08 3.48 ;
        RECT  4.82 2.29 5.10 2.57 ;
        RECT  4.88 2.29 5.04 3.48 ;
        RECT  3.66 1.84 3.94 2.12 ;
        RECT  3.72 1.84 3.88 3.48 ;
        RECT  1.66 2.29 1.94 2.57 ;
        RECT  1.72 2.29 1.88 3.48 ;
        RECT  0.62 2.29 0.90 2.57 ;
        RECT  0.68 2.29 0.84 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.08 0.75 0.58 1.03 ;
        RECT  2.44 1.40 2.88 1.68 ;
        RECT  0.08 0.75 0.24 2.13 ;
        RECT  2.44 1.40 2.60 2.13 ;
        RECT  0.08 1.97 2.60 2.13 ;
        RECT  0.16 1.97 0.32 2.57 ;
        RECT  1.20 1.97 1.36 2.57 ;
        RECT  2.24 1.97 2.40 2.57 ;
        RECT  0.10 2.29 0.38 2.57 ;
        RECT  1.14 2.29 1.42 2.57 ;
        RECT  2.18 2.29 2.46 2.57 ;
        RECT  3.20 0.96 3.56 1.24 ;
        RECT  3.20 1.46 4.28 1.62 ;
        RECT  4.00 1.40 4.28 1.68 ;
        RECT  3.20 0.96 3.36 2.00 ;
        RECT  2.76 1.84 3.36 2.00 ;
        RECT  2.76 1.84 3.04 2.12 ;
        RECT  4.46 0.44 4.74 0.72 ;
        RECT  4.46 0.56 5.32 0.72 ;
        RECT  5.04 0.56 5.32 0.91 ;
        RECT  5.10 0.56 5.26 1.23 ;
        RECT  5.10 1.07 6.74 1.23 ;
        RECT  6.58 1.07 6.74 2.13 ;
        RECT  5.46 1.97 6.74 2.13 ;
        RECT  6.50 1.97 6.66 2.57 ;
        RECT  5.46 1.97 5.62 2.57 ;
        RECT  5.34 2.29 5.62 2.57 ;
        RECT  6.38 2.29 6.66 2.57 ;
    END
END NAND8SP1V1_0

MACRO NAND6SP8V1_0
    CLASS CORE ;
    FOREIGN NAND6SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN6
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.64 1.39 7.92 1.81 ;
        RECT  7.56 1.46 7.92 1.74 ;
        END
    END IN6
    PIN IN5
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.92 1.39 7.20 1.81 ;
        END
    END IN5
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.46 1.39 6.74 1.81 ;
        RECT  6.44 1.46 6.74 1.74 ;
        END
    END IN4
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.39 0.68 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.88 1.39 1.16 1.81 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.32 1.46 1.74 1.74 ;
        END
    END IN3
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 14.93  LAYER ME1  ;
        ANTENNADIFFAREA 7.98  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.89  LAYER ME1  ;
        ANTENNAMAXAREACAR 16.73  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.85 0.66 5.14 1.24 ;
        RECT  4.72 1.84 5.01 2.42 ;
        RECT  4.85 0.66 5.01 2.42 ;
        RECT  3.92 1.52 5.01 1.68 ;
        RECT  3.82 0.66 4.10 1.24 ;
        RECT  3.92 0.66 4.08 2.00 ;
        RECT  3.68 1.84 3.96 2.42 ;
        END
    END OUT
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 8.00 0.28 ;
        RECT  7.54 -0.28 7.82 0.32 ;
        RECT  7.48 0.63 7.76 0.91 ;
        RECT  7.54 -0.28 7.70 0.91 ;
        RECT  5.38 0.66 5.66 1.24 ;
        RECT  5.40 -0.28 5.56 1.24 ;
        RECT  4.34 0.66 4.62 1.24 ;
        RECT  4.36 -0.28 4.52 1.24 ;
        RECT  3.26 0.54 3.54 1.24 ;
        RECT  3.28 -0.28 3.44 1.24 ;
        RECT  2.22 0.54 2.50 1.24 ;
        RECT  2.28 -0.28 2.44 1.24 ;
        RECT  1.52 0.85 1.80 1.13 ;
        RECT  1.58 -0.28 1.74 1.13 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 8.00 3.48 ;
        RECT  7.54 2.88 7.82 3.48 ;
        RECT  7.10 2.29 7.38 2.57 ;
        RECT  7.16 2.29 7.32 3.48 ;
        RECT  6.06 2.29 6.34 2.57 ;
        RECT  6.12 2.29 6.28 3.48 ;
        RECT  5.24 2.14 5.52 2.42 ;
        RECT  5.30 2.14 5.46 3.48 ;
        RECT  4.20 2.14 4.48 2.42 ;
        RECT  4.26 2.14 4.42 3.48 ;
        RECT  3.12 1.84 3.40 2.54 ;
        RECT  3.18 1.84 3.34 3.48 ;
        RECT  1.66 2.29 1.94 2.57 ;
        RECT  1.72 2.29 1.88 3.48 ;
        RECT  0.62 2.29 0.90 2.57 ;
        RECT  0.68 2.29 0.84 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.08 0.85 0.52 1.13 ;
        RECT  1.90 1.40 2.34 1.68 ;
        RECT  0.08 0.85 0.24 2.13 ;
        RECT  1.90 1.40 2.06 2.13 ;
        RECT  0.08 1.97 2.06 2.13 ;
        RECT  0.16 1.97 0.32 2.57 ;
        RECT  1.14 1.97 1.30 2.57 ;
        RECT  0.10 2.29 0.38 2.57 ;
        RECT  1.14 2.29 1.42 2.57 ;
        RECT  2.66 0.54 3.02 1.24 ;
        RECT  2.66 1.46 3.76 1.62 ;
        RECT  3.48 1.40 3.76 1.68 ;
        RECT  2.66 0.54 2.82 2.00 ;
        RECT  2.22 1.84 2.82 2.00 ;
        RECT  2.22 1.84 2.50 2.54 ;
        RECT  5.96 0.63 6.48 0.91 ;
        RECT  5.96 0.63 6.12 2.13 ;
        RECT  5.68 1.85 6.12 2.13 ;
        RECT  5.68 1.97 7.78 2.13 ;
        RECT  7.62 1.97 7.78 2.57 ;
        RECT  6.70 1.97 6.86 2.57 ;
        RECT  6.58 2.29 6.86 2.57 ;
        RECT  7.62 2.29 7.90 2.57 ;
    END
END NAND6SP8V1_0

MACRO NAND6SP4V1_0
    CLASS CORE ;
    FOREIGN NAND6SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN5
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.66 1.39 5.94 1.81 ;
        END
    END IN5
    PIN IN6
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.44 1.39 6.72 1.81 ;
        RECT  6.26 1.46 6.72 1.74 ;
        END
    END IN6
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.22 1.39 5.50 1.81 ;
        RECT  5.14 1.46 5.50 1.74 ;
        END
    END IN4
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 12.01  LAYER ME1  ;
        ANTENNADIFFAREA 6.14  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.56  LAYER ME1  ;
        ANTENNAMAXAREACAR 21.57  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.90 1.52 4.28 1.68 ;
        RECT  3.90 0.66 4.06 2.00 ;
        RECT  3.64 1.84 3.92 2.42 ;
        RECT  3.78 0.66 4.06 1.24 ;
        END
    END OUT
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.32 1.46 1.74 1.74 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.88 1.39 1.16 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.39 0.68 1.81 ;
        END
    END IN1
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 6.80 3.48 ;
        RECT  6.34 2.88 6.62 3.48 ;
        RECT  5.80 2.29 6.08 2.57 ;
        RECT  5.86 2.29 6.02 3.48 ;
        RECT  4.76 2.29 5.04 2.57 ;
        RECT  4.82 2.29 4.98 3.48 ;
        RECT  4.16 2.14 4.44 2.42 ;
        RECT  4.22 2.14 4.38 3.48 ;
        RECT  3.12 1.84 3.40 2.42 ;
        RECT  3.18 1.84 3.34 3.48 ;
        RECT  1.66 2.29 1.94 2.57 ;
        RECT  1.72 2.29 1.88 3.48 ;
        RECT  0.62 2.29 0.90 2.57 ;
        RECT  0.68 2.29 0.84 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 6.80 0.28 ;
        RECT  6.24 -0.28 6.62 0.32 ;
        RECT  6.18 0.63 6.46 0.91 ;
        RECT  6.24 -0.28 6.40 0.91 ;
        RECT  4.30 0.66 4.58 1.24 ;
        RECT  4.36 -0.28 4.52 1.24 ;
        RECT  3.26 0.66 3.54 1.24 ;
        RECT  3.32 -0.28 3.48 1.24 ;
        RECT  2.22 0.66 2.50 1.24 ;
        RECT  2.28 -0.28 2.44 1.24 ;
        RECT  1.52 0.85 1.80 1.13 ;
        RECT  1.58 -0.28 1.74 1.13 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.08 0.85 0.52 1.13 ;
        RECT  1.90 1.40 2.34 1.68 ;
        RECT  0.08 0.85 0.24 2.13 ;
        RECT  1.90 1.40 2.06 2.13 ;
        RECT  0.08 1.97 2.06 2.13 ;
        RECT  0.16 1.97 0.32 2.57 ;
        RECT  1.14 1.97 1.30 2.57 ;
        RECT  0.10 2.29 0.38 2.57 ;
        RECT  1.14 2.29 1.42 2.57 ;
        RECT  2.66 0.66 3.02 1.24 ;
        RECT  2.66 1.46 3.74 1.62 ;
        RECT  3.46 1.40 3.74 1.68 ;
        RECT  2.66 0.66 2.82 2.00 ;
        RECT  2.22 1.84 2.82 2.00 ;
        RECT  2.22 1.84 2.50 2.42 ;
        RECT  4.80 0.63 5.18 0.91 ;
        RECT  4.80 0.63 4.96 2.13 ;
        RECT  4.60 1.85 4.96 2.13 ;
        RECT  4.60 1.97 6.48 2.13 ;
        RECT  6.32 1.97 6.48 2.57 ;
        RECT  5.40 1.97 5.56 2.57 ;
        RECT  5.28 2.29 5.56 2.57 ;
        RECT  6.32 2.29 6.60 2.57 ;
    END
END NAND6SP4V1_0

MACRO NAND6SP2V1_0
    CLASS CORE ;
    FOREIGN NAND6SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN6
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.04 1.39 6.32 1.81 ;
        RECT  6.02 1.46 6.32 1.74 ;
        END
    END IN6
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.39 0.68 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.88 1.39 1.16 1.81 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.32 1.46 1.74 1.74 ;
        END
    END IN3
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.82 1.39 5.10 1.81 ;
        END
    END IN4
    PIN IN5
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.30 1.39 5.58 1.81 ;
        END
    END IN5
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 11.08  LAYER ME1  ;
        ANTENNADIFFAREA 5.18  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.34  LAYER ME1  ;
        ANTENNAMAXAREACAR 32.97  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.94 1.52 4.28 1.68 ;
        RECT  3.94 0.64 4.10 2.00 ;
        RECT  3.68 1.84 3.96 2.12 ;
        RECT  3.82 0.64 4.10 1.24 ;
        END
    END OUT
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 6.40 0.28 ;
        RECT  5.94 -0.28 6.22 0.32 ;
        RECT  5.88 0.63 6.16 0.91 ;
        RECT  5.94 -0.28 6.10 0.91 ;
        RECT  3.30 0.64 3.58 1.24 ;
        RECT  3.36 -0.28 3.52 1.24 ;
        RECT  2.22 0.84 2.50 1.24 ;
        RECT  2.28 -0.28 2.44 1.24 ;
        RECT  1.52 0.85 1.80 1.13 ;
        RECT  1.58 -0.28 1.74 1.13 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 6.40 3.48 ;
        RECT  5.94 2.88 6.22 3.48 ;
        RECT  5.50 2.29 5.78 2.57 ;
        RECT  5.56 2.29 5.72 3.48 ;
        RECT  4.42 2.62 4.70 3.48 ;
        RECT  3.16 1.84 3.44 2.44 ;
        RECT  3.18 1.84 3.34 3.48 ;
        RECT  1.66 2.29 1.94 2.57 ;
        RECT  1.72 2.29 1.88 3.48 ;
        RECT  0.62 2.29 0.90 2.57 ;
        RECT  0.68 2.29 0.84 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.08 0.85 0.52 1.13 ;
        RECT  1.90 1.40 2.34 1.68 ;
        RECT  0.08 0.85 0.24 2.13 ;
        RECT  1.90 1.40 2.06 2.13 ;
        RECT  0.08 1.97 2.06 2.13 ;
        RECT  0.16 1.97 0.32 2.57 ;
        RECT  1.14 1.97 1.30 2.57 ;
        RECT  0.10 2.29 0.38 2.57 ;
        RECT  1.14 2.29 1.42 2.57 ;
        RECT  2.66 0.84 3.02 1.24 ;
        RECT  2.66 1.46 3.77 1.62 ;
        RECT  3.49 1.40 3.77 1.68 ;
        RECT  2.66 0.84 2.82 2.00 ;
        RECT  2.22 1.84 2.82 2.00 ;
        RECT  2.22 1.84 2.50 2.24 ;
        RECT  4.50 0.63 4.88 0.91 ;
        RECT  4.50 0.63 4.66 2.13 ;
        RECT  4.44 1.97 6.18 2.13 ;
        RECT  4.44 1.97 4.60 2.43 ;
        RECT  6.02 1.97 6.18 2.57 ;
        RECT  4.16 2.15 4.60 2.43 ;
        RECT  5.10 1.97 5.26 2.57 ;
        RECT  4.98 2.29 5.26 2.57 ;
        RECT  6.02 2.29 6.30 2.57 ;
    END
END NAND6SP2V1_0

MACRO NAND6SP1V1_0
    CLASS CORE ;
    FOREIGN NAND6SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 11.13  LAYER ME1  ;
        ANTENNADIFFAREA 4.47  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        ANTENNAMAXAREACAR 55.19  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.64 1.84 4.28 2.00 ;
        RECT  4.12 1.08 4.28 2.00 ;
        RECT  3.78 1.08 4.28 1.24 ;
        RECT  3.78 0.96 4.06 1.24 ;
        RECT  3.64 1.84 3.92 2.12 ;
        END
    END OUT
    PIN IN5
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.18 1.39 5.50 1.81 ;
        END
    END IN5
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.46 1.39 4.74 1.81 ;
        END
    END IN4
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.32 1.46 1.74 1.74 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.88 1.39 1.16 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.39 0.68 1.81 ;
        END
    END IN1
    PIN IN6
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.66 1.39 5.94 1.81 ;
        END
    END IN6
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 6.40 3.48 ;
        RECT  5.94 2.88 6.22 3.48 ;
        RECT  5.32 2.29 5.60 2.57 ;
        RECT  5.38 2.29 5.54 3.48 ;
        RECT  4.28 2.29 4.56 2.57 ;
        RECT  4.34 2.29 4.50 3.48 ;
        RECT  3.12 1.84 3.40 2.12 ;
        RECT  3.18 1.84 3.34 3.48 ;
        RECT  1.66 2.29 1.94 2.57 ;
        RECT  1.72 2.29 1.88 3.48 ;
        RECT  0.62 2.29 0.90 2.57 ;
        RECT  0.68 2.29 0.84 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 6.40 0.28 ;
        RECT  5.76 -0.28 6.22 0.32 ;
        RECT  5.70 0.63 5.98 0.91 ;
        RECT  5.76 -0.28 5.92 0.91 ;
        RECT  3.26 0.96 3.54 1.24 ;
        RECT  3.32 -0.28 3.48 1.24 ;
        RECT  2.22 0.96 2.50 1.24 ;
        RECT  2.28 -0.28 2.44 1.24 ;
        RECT  1.52 0.85 1.80 1.13 ;
        RECT  1.58 -0.28 1.74 1.13 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.08 0.85 0.52 1.13 ;
        RECT  1.90 1.40 2.34 1.68 ;
        RECT  0.08 0.85 0.24 2.13 ;
        RECT  1.90 1.40 2.06 2.13 ;
        RECT  0.08 1.97 2.06 2.13 ;
        RECT  0.16 1.97 0.32 2.57 ;
        RECT  1.14 1.97 1.30 2.57 ;
        RECT  0.10 2.29 0.38 2.57 ;
        RECT  1.14 2.29 1.42 2.57 ;
        RECT  2.66 0.96 3.02 1.24 ;
        RECT  2.66 1.46 3.74 1.62 ;
        RECT  3.46 1.40 3.74 1.68 ;
        RECT  2.66 0.96 2.82 2.00 ;
        RECT  2.22 1.84 2.82 2.00 ;
        RECT  2.22 1.84 2.50 2.12 ;
        RECT  3.92 0.44 4.20 0.72 ;
        RECT  3.92 0.56 4.70 0.72 ;
        RECT  4.42 0.56 4.70 0.91 ;
        RECT  4.54 0.56 4.70 1.23 ;
        RECT  4.54 1.07 6.26 1.23 ;
        RECT  6.10 1.07 6.26 2.13 ;
        RECT  4.92 1.97 6.26 2.13 ;
        RECT  5.96 1.97 6.12 2.57 ;
        RECT  4.92 1.97 5.08 2.57 ;
        RECT  4.80 2.29 5.08 2.57 ;
        RECT  5.84 2.29 6.12 2.57 ;
    END
END NAND6SP1V1_0

MACRO NAND5SP8V1_0
    CLASS CORE ;
    FOREIGN NAND5SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.06 1.39 6.34 1.81 ;
        END
    END IN4
    PIN IN5
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.86 1.39 7.14 1.81 ;
        END
    END IN5
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 14.23  LAYER ME1  ;
        ANTENNADIFFAREA 7.92  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.89  LAYER ME1  ;
        ANTENNAMAXAREACAR 15.94  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.85 0.64 5.14 1.22 ;
        RECT  4.72 1.84 5.01 2.42 ;
        RECT  4.85 0.64 5.01 2.42 ;
        RECT  3.94 1.52 5.01 1.68 ;
        RECT  3.94 0.64 4.10 2.00 ;
        RECT  3.68 1.84 3.96 2.42 ;
        RECT  3.82 0.64 4.10 1.22 ;
        END
    END OUT
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.32 1.46 1.74 1.74 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.88 1.39 1.16 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.39 0.68 1.81 ;
        END
    END IN1
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 7.60 3.48 ;
        RECT  7.10 2.88 7.42 3.48 ;
        RECT  7.04 1.97 7.32 2.25 ;
        RECT  7.10 1.97 7.26 3.48 ;
        RECT  6.00 2.62 6.28 3.48 ;
        RECT  5.24 1.84 5.52 2.42 ;
        RECT  5.30 1.84 5.46 3.48 ;
        RECT  4.20 2.14 4.48 2.42 ;
        RECT  4.26 2.14 4.42 3.48 ;
        RECT  3.12 1.84 3.40 2.54 ;
        RECT  3.18 1.84 3.34 3.48 ;
        RECT  1.66 2.29 1.94 2.57 ;
        RECT  1.72 2.29 1.88 3.48 ;
        RECT  0.62 2.29 0.90 2.57 ;
        RECT  0.68 2.29 0.84 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 7.60 0.28 ;
        RECT  7.03 -0.28 7.42 0.32 ;
        RECT  6.97 0.95 7.25 1.23 ;
        RECT  7.03 -0.28 7.19 1.23 ;
        RECT  5.38 0.64 5.66 1.22 ;
        RECT  5.44 -0.28 5.60 1.22 ;
        RECT  4.34 0.64 4.62 1.22 ;
        RECT  4.40 -0.28 4.56 1.22 ;
        RECT  3.26 0.52 3.54 1.22 ;
        RECT  3.32 -0.28 3.48 1.22 ;
        RECT  2.22 0.52 2.50 1.22 ;
        RECT  2.28 -0.28 2.44 1.22 ;
        RECT  1.52 0.85 1.80 1.13 ;
        RECT  1.58 -0.28 1.74 1.13 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.08 0.85 0.52 1.13 ;
        RECT  1.90 1.40 2.34 1.68 ;
        RECT  0.08 0.85 0.24 2.13 ;
        RECT  1.90 1.40 2.06 2.13 ;
        RECT  0.08 1.97 2.06 2.13 ;
        RECT  0.16 1.97 0.32 2.57 ;
        RECT  1.14 1.97 1.30 2.57 ;
        RECT  0.10 2.29 0.38 2.57 ;
        RECT  1.14 2.29 1.42 2.57 ;
        RECT  2.74 0.52 3.02 1.22 ;
        RECT  2.66 1.46 3.76 1.62 ;
        RECT  3.48 1.40 3.76 1.68 ;
        RECT  2.66 0.66 2.82 2.00 ;
        RECT  2.22 1.84 2.82 2.00 ;
        RECT  2.22 1.84 2.50 2.54 ;
        RECT  6.07 0.95 6.35 1.23 ;
        RECT  6.07 1.07 6.66 1.23 ;
        RECT  6.50 1.07 6.66 2.32 ;
        RECT  6.50 1.97 6.80 2.32 ;
        RECT  5.68 2.16 6.80 2.32 ;
        RECT  5.68 2.16 5.96 2.44 ;
    END
END NAND5SP8V1_0

MACRO NAND5SP4V1_0
    CLASS CORE ;
    FOREIGN NAND5SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.39 0.68 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.88 1.39 1.16 1.81 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.32 1.46 1.74 1.74 ;
        END
    END IN3
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.86 1.39 5.14 1.81 ;
        END
    END IN4
    PIN IN5
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.69 1.39 5.97 1.81 ;
        END
    END IN5
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 11.32  LAYER ME1  ;
        ANTENNADIFFAREA 6.21  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER ME1  ;
        ANTENNAMAXAREACAR 19.99  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.94 1.52 4.28 1.68 ;
        RECT  3.94 0.64 4.10 2.00 ;
        RECT  3.68 1.84 3.96 2.44 ;
        RECT  3.82 0.64 4.10 1.24 ;
        END
    END OUT
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 6.40 0.28 ;
        RECT  5.94 -0.28 6.22 0.32 ;
        RECT  5.93 0.95 6.21 1.23 ;
        RECT  5.99 -0.28 6.15 1.23 ;
        RECT  4.34 0.64 4.62 1.24 ;
        RECT  4.40 -0.28 4.56 1.24 ;
        RECT  3.30 0.64 3.58 1.24 ;
        RECT  3.36 -0.28 3.52 1.24 ;
        RECT  2.22 0.66 2.50 1.24 ;
        RECT  2.28 -0.28 2.44 1.24 ;
        RECT  1.52 0.85 1.80 1.13 ;
        RECT  1.58 -0.28 1.74 1.13 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 6.40 3.48 ;
        RECT  6.00 1.97 6.28 2.25 ;
        RECT  5.94 2.88 6.22 3.48 ;
        RECT  6.06 1.97 6.22 3.48 ;
        RECT  4.96 2.62 5.24 3.48 ;
        RECT  4.20 2.16 4.48 2.44 ;
        RECT  4.26 2.16 4.42 3.48 ;
        RECT  3.16 1.84 3.44 2.44 ;
        RECT  3.22 1.84 3.38 3.48 ;
        RECT  1.66 2.29 1.94 2.57 ;
        RECT  1.72 2.29 1.88 3.48 ;
        RECT  0.62 2.29 0.90 2.57 ;
        RECT  0.68 2.29 0.84 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.08 0.85 0.52 1.13 ;
        RECT  1.90 1.40 2.34 1.68 ;
        RECT  0.08 0.85 0.24 2.13 ;
        RECT  1.90 1.40 2.06 2.13 ;
        RECT  0.08 1.97 2.06 2.13 ;
        RECT  0.16 1.97 0.32 2.57 ;
        RECT  1.14 1.97 1.30 2.57 ;
        RECT  0.10 2.29 0.38 2.57 ;
        RECT  1.14 2.29 1.42 2.57 ;
        RECT  2.66 0.66 3.02 1.24 ;
        RECT  2.66 1.46 3.76 1.62 ;
        RECT  3.48 1.40 3.76 1.68 ;
        RECT  2.66 0.66 2.82 2.00 ;
        RECT  2.22 1.84 2.82 2.00 ;
        RECT  2.22 1.84 2.50 2.42 ;
        RECT  5.03 0.95 5.31 1.23 ;
        RECT  5.03 1.07 5.48 1.23 ;
        RECT  5.32 1.07 5.48 2.32 ;
        RECT  5.32 1.97 5.76 2.32 ;
        RECT  4.64 2.16 5.76 2.32 ;
        RECT  4.64 2.16 4.92 2.44 ;
    END
END NAND5SP4V1_0

MACRO NAND5SP2V1_0
    CLASS CORE ;
    FOREIGN NAND5SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 10.35  LAYER ME1  ;
        ANTENNADIFFAREA 5.06  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.34  LAYER ME1  ;
        ANTENNAMAXAREACAR 30.82  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.68 1.84 4.28 2.00 ;
        RECT  4.12 1.08 4.28 2.00 ;
        RECT  3.82 1.08 4.28 1.24 ;
        RECT  3.82 0.64 4.10 1.24 ;
        RECT  3.68 1.84 3.96 2.44 ;
        END
    END OUT
    PIN IN5
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.26 1.39 5.54 1.81 ;
        END
    END IN5
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.46 1.39 4.74 1.81 ;
        END
    END IN4
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.32 1.46 1.74 1.74 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.88 1.39 1.16 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.39 0.68 1.81 ;
        END
    END IN1
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 6.00 3.48 ;
        RECT  5.54 2.88 5.82 3.48 ;
        RECT  5.48 1.97 5.76 2.25 ;
        RECT  5.54 1.97 5.70 3.48 ;
        RECT  4.44 2.62 4.72 3.48 ;
        RECT  3.16 1.84 3.44 2.44 ;
        RECT  3.22 1.84 3.38 3.48 ;
        RECT  1.66 2.29 1.94 2.57 ;
        RECT  1.72 2.29 1.88 3.48 ;
        RECT  0.62 2.29 0.90 2.57 ;
        RECT  0.68 2.29 0.84 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 6.00 0.28 ;
        RECT  5.47 -0.28 5.82 0.32 ;
        RECT  5.41 0.95 5.69 1.23 ;
        RECT  5.47 -0.28 5.63 1.23 ;
        RECT  3.30 0.64 3.58 1.24 ;
        RECT  3.36 -0.28 3.52 1.24 ;
        RECT  2.22 0.84 2.50 1.24 ;
        RECT  2.28 -0.28 2.44 1.24 ;
        RECT  1.52 0.85 1.80 1.13 ;
        RECT  1.58 -0.28 1.74 1.13 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.08 0.85 0.52 1.13 ;
        RECT  1.90 1.40 2.34 1.68 ;
        RECT  0.08 0.85 0.24 2.13 ;
        RECT  1.90 1.40 2.06 2.13 ;
        RECT  0.08 1.97 2.06 2.13 ;
        RECT  0.16 1.97 0.32 2.57 ;
        RECT  1.14 1.97 1.30 2.57 ;
        RECT  0.10 2.29 0.38 2.57 ;
        RECT  1.14 2.29 1.42 2.57 ;
        RECT  2.66 0.84 3.02 1.24 ;
        RECT  2.66 1.46 3.76 1.62 ;
        RECT  3.48 1.40 3.76 1.68 ;
        RECT  2.66 0.84 2.82 2.00 ;
        RECT  2.22 1.84 2.82 2.00 ;
        RECT  2.22 1.84 2.50 2.24 ;
        RECT  4.51 0.95 4.79 1.23 ;
        RECT  4.51 1.07 5.06 1.23 ;
        RECT  4.90 1.07 5.06 2.32 ;
        RECT  4.90 1.97 5.24 2.32 ;
        RECT  4.12 2.16 5.24 2.32 ;
        RECT  4.12 2.16 4.40 2.44 ;
    END
END NAND5SP2V1_0

MACRO NAND5SP1V1_0
    CLASS CORE ;
    FOREIGN NAND5SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.39 0.68 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.88 1.39 1.16 1.81 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.32 1.46 1.74 1.74 ;
        END
    END IN3
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.46 1.39 4.74 1.81 ;
        END
    END IN4
    PIN IN5
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.26 1.39 5.54 1.81 ;
        END
    END IN5
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 10.22  LAYER ME1  ;
        ANTENNADIFFAREA 4.16  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        ANTENNAMAXAREACAR 50.70  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.64 1.84 4.28 2.00 ;
        RECT  4.12 1.08 4.28 2.00 ;
        RECT  3.78 1.08 4.28 1.24 ;
        RECT  3.78 0.96 4.06 1.24 ;
        RECT  3.64 1.84 3.92 2.12 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 6.00 3.48 ;
        RECT  5.38 2.88 5.82 3.48 ;
        RECT  5.32 2.16 5.60 2.44 ;
        RECT  5.38 2.16 5.54 3.48 ;
        RECT  4.28 2.16 4.56 2.44 ;
        RECT  4.34 2.16 4.50 3.48 ;
        RECT  3.12 1.84 3.40 2.12 ;
        RECT  3.18 1.84 3.34 3.48 ;
        RECT  1.66 2.29 1.94 2.57 ;
        RECT  1.72 2.29 1.88 3.48 ;
        RECT  0.62 2.29 0.90 2.57 ;
        RECT  0.68 2.29 0.84 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 6.00 0.28 ;
        RECT  5.31 -0.28 5.82 0.32 ;
        RECT  5.25 0.65 5.53 0.93 ;
        RECT  5.31 -0.28 5.47 0.93 ;
        RECT  3.26 0.96 3.54 1.24 ;
        RECT  3.32 -0.28 3.48 1.24 ;
        RECT  2.22 0.96 2.50 1.24 ;
        RECT  2.28 -0.28 2.44 1.24 ;
        RECT  1.52 0.85 1.80 1.13 ;
        RECT  1.58 -0.28 1.74 1.13 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.08 0.85 0.52 1.13 ;
        RECT  1.90 1.40 2.34 1.68 ;
        RECT  0.08 0.85 0.24 2.13 ;
        RECT  1.90 1.40 2.06 2.13 ;
        RECT  0.08 1.97 2.06 2.13 ;
        RECT  0.16 1.97 0.32 2.57 ;
        RECT  1.14 1.97 1.30 2.57 ;
        RECT  0.10 2.29 0.38 2.57 ;
        RECT  1.14 2.29 1.42 2.57 ;
        RECT  2.66 0.96 3.02 1.24 ;
        RECT  2.66 1.46 3.74 1.62 ;
        RECT  3.46 1.40 3.74 1.68 ;
        RECT  2.66 0.96 2.82 2.00 ;
        RECT  2.22 1.84 2.82 2.00 ;
        RECT  2.22 1.84 2.50 2.12 ;
        RECT  3.92 0.44 4.20 0.72 ;
        RECT  3.92 0.56 4.63 0.72 ;
        RECT  4.35 0.56 4.63 0.93 ;
        RECT  4.35 0.77 5.06 0.93 ;
        RECT  4.90 0.77 5.06 2.44 ;
        RECT  4.80 2.16 5.08 2.44 ;
    END
END NAND5SP1V1_0

MACRO NAND4SP9V1_0
    CLASS CORE ;
    FOREIGN NAND4SP9V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.43 0.38 1.85 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.88 1.43 1.16 1.85 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.32 1.43 1.64 1.85 ;
        END
    END IN3
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.12 1.76 2.40 2.18 ;
        END
    END IN4
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 7.40  LAYER ME1  ;
        ANTENNADIFFAREA 3.82  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.27  LAYER ME1  ;
        ANTENNAMAXAREACAR 27.05  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.78 1.84 4.28 2.12 ;
        RECT  4.12 0.96 4.28 2.12 ;
        RECT  3.78 0.96 4.28 1.24 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.40 3.48 ;
        RECT  3.94 2.88 4.22 3.48 ;
        RECT  3.26 2.26 3.54 2.54 ;
        RECT  3.32 2.26 3.48 3.48 ;
        RECT  2.18 2.34 2.46 2.62 ;
        RECT  2.24 2.34 2.40 3.48 ;
        RECT  1.14 2.34 1.42 2.62 ;
        RECT  1.20 2.34 1.36 3.48 ;
        RECT  0.10 2.34 0.38 2.62 ;
        RECT  0.16 2.34 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.40 0.28 ;
        RECT  3.94 -0.28 4.22 0.32 ;
        RECT  3.26 0.54 3.54 0.82 ;
        RECT  3.32 -0.28 3.48 0.82 ;
        RECT  1.97 0.66 2.25 0.94 ;
        RECT  2.03 -0.28 2.19 0.94 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.31 0.66 0.59 0.94 ;
        RECT  0.43 0.66 0.59 1.27 ;
        RECT  0.43 1.11 1.96 1.27 ;
        RECT  1.80 1.44 3.20 1.60 ;
        RECT  2.92 1.40 3.20 1.68 ;
        RECT  1.80 1.11 1.96 2.18 ;
        RECT  0.74 2.02 1.96 2.18 ;
        RECT  1.66 2.02 1.82 2.62 ;
        RECT  0.74 2.02 0.90 2.62 ;
        RECT  0.62 2.34 0.90 2.62 ;
        RECT  1.66 2.34 1.94 2.62 ;
        RECT  2.70 0.70 2.98 0.98 ;
        RECT  2.82 0.70 2.98 1.24 ;
        RECT  2.82 1.08 3.60 1.24 ;
        RECT  3.44 1.40 3.72 1.68 ;
        RECT  3.44 1.08 3.60 2.00 ;
        RECT  2.82 1.84 3.60 2.00 ;
        RECT  2.82 1.84 2.98 2.38 ;
        RECT  2.70 2.10 2.98 2.38 ;
    END
END NAND4SP9V1_0

MACRO NAND4SP8V1_0
    CLASS CORE ;
    FOREIGN NAND4SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.58  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.28 1.39 1.56 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.58  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.86 1.39 3.14 1.81 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.58  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.46 1.39 4.74 1.81 ;
        END
    END IN3
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.46  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.99 1.44 6.41 1.72 ;
        END
    END IN4
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 12.13  LAYER ME1  ;
        ANTENNADIFFAREA 10.44  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.86 2.10 6.14 2.38 ;
        RECT  5.86 1.88 6.02 2.38 ;
        RECT  4.90 1.88 6.02 2.04 ;
        RECT  4.78 2.04 5.06 2.38 ;
        RECT  0.52 2.04 5.06 2.20 ;
        RECT  3.74 2.04 4.02 2.38 ;
        RECT  2.70 2.04 2.98 2.38 ;
        RECT  1.66 2.04 1.94 2.38 ;
        RECT  0.10 0.88 1.42 1.04 ;
        RECT  1.14 0.76 1.42 1.04 ;
        RECT  0.62 2.04 0.90 2.38 ;
        RECT  0.52 0.88 0.68 2.20 ;
        RECT  0.10 0.76 0.38 1.04 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 6.80 3.48 ;
        RECT  6.38 2.20 6.66 2.48 ;
        RECT  6.34 2.88 6.62 3.48 ;
        RECT  6.44 2.20 6.60 3.48 ;
        RECT  5.34 2.20 5.62 2.48 ;
        RECT  5.40 2.20 5.56 3.48 ;
        RECT  4.26 2.36 4.54 2.64 ;
        RECT  4.32 2.36 4.48 3.48 ;
        RECT  3.22 2.36 3.50 2.64 ;
        RECT  3.28 2.36 3.44 3.48 ;
        RECT  2.18 2.36 2.46 2.64 ;
        RECT  2.24 2.36 2.40 3.48 ;
        RECT  1.14 2.36 1.42 2.64 ;
        RECT  1.20 2.36 1.36 3.48 ;
        RECT  0.10 2.36 0.38 2.64 ;
        RECT  0.16 2.36 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 6.80 0.28 ;
        RECT  6.38 0.60 6.66 0.88 ;
        RECT  6.34 -0.28 6.62 0.32 ;
        RECT  6.44 -0.28 6.60 0.88 ;
        RECT  5.34 0.60 5.62 0.88 ;
        RECT  5.40 -0.28 5.56 0.88 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.44 1.94 0.60 ;
        RECT  0.62 0.44 0.90 0.72 ;
        RECT  1.66 0.44 1.94 0.72 ;
        RECT  1.78 0.44 1.94 1.04 ;
        RECT  2.70 0.76 2.98 1.04 ;
        RECT  1.78 0.88 2.98 1.04 ;
        RECT  2.18 0.44 3.50 0.60 ;
        RECT  2.18 0.44 2.46 0.72 ;
        RECT  3.22 0.44 3.50 0.72 ;
        RECT  3.34 0.44 3.50 1.04 ;
        RECT  4.26 0.76 4.54 1.04 ;
        RECT  3.34 0.88 4.54 1.04 ;
        RECT  3.74 0.44 5.06 0.60 ;
        RECT  3.74 0.44 4.02 0.72 ;
        RECT  4.78 0.44 5.06 0.72 ;
        RECT  4.90 0.44 5.06 1.20 ;
        RECT  5.86 0.76 6.14 1.04 ;
        RECT  4.90 1.04 6.02 1.20 ;
    END
END NAND4SP8V1_0

MACRO NAND4SP2V1_0
    CLASS CORE ;
    FOREIGN NAND4SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 2.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.14  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.34 0.68 1.76 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.14  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.88 1.34 1.16 1.76 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.14  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.37 1.38 1.65 1.80 ;
        RECT  1.32 1.52 1.65 1.68 ;
        END
    END IN3
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.14  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.00 1.34 2.28 1.76 ;
        END
    END IN4
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 3.63  LAYER ME1  ;
        ANTENNADIFFAREA 3.27  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.66 2.38 1.94 2.66 ;
        RECT  1.66 2.06 1.82 2.66 ;
        RECT  0.74 2.06 1.82 2.22 ;
        RECT  0.62 2.38 0.90 2.66 ;
        RECT  0.74 1.92 0.90 2.66 ;
        RECT  0.08 1.92 0.90 2.08 ;
        RECT  0.08 0.82 0.50 1.10 ;
        RECT  0.08 0.82 0.24 2.08 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 2.80 3.48 ;
        RECT  2.24 2.88 2.62 3.48 ;
        RECT  2.18 2.38 2.46 2.66 ;
        RECT  2.24 2.38 2.40 3.48 ;
        RECT  1.14 2.38 1.42 2.66 ;
        RECT  1.20 2.38 1.36 3.48 ;
        RECT  0.10 2.38 0.38 2.66 ;
        RECT  0.16 2.38 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 2.80 0.28 ;
        RECT  2.34 -0.28 2.62 0.32 ;
        RECT  1.88 0.50 2.16 0.78 ;
        RECT  1.95 -0.28 2.11 0.78 ;
        END
    END GND!
END NAND4SP2V1_0

MACRO NAND4SP1V1_0
    CLASS CORE ;
    FOREIGN NAND4SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 2.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.26 0.68 1.68 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.88 1.26 1.16 1.68 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.32 1.40 1.74 1.68 ;
        END
    END IN3
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.06 1.26 2.34 1.68 ;
        END
    END IN4
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 3.72  LAYER ME1  ;
        ANTENNADIFFAREA 1.97  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.66 2.24 1.94 2.52 ;
        RECT  0.08 1.92 1.88 2.08 ;
        RECT  1.66 1.92 1.82 2.52 ;
        RECT  0.62 2.24 0.90 2.52 ;
        RECT  0.74 1.92 0.90 2.52 ;
        RECT  0.08 0.78 0.59 0.94 ;
        RECT  0.31 0.66 0.59 0.94 ;
        RECT  0.08 0.78 0.24 2.08 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 2.80 3.48 ;
        RECT  2.24 2.88 2.62 3.48 ;
        RECT  2.18 2.24 2.46 2.52 ;
        RECT  2.24 2.24 2.40 3.48 ;
        RECT  1.14 2.24 1.42 2.52 ;
        RECT  1.20 2.24 1.36 3.48 ;
        RECT  0.10 2.24 0.38 2.52 ;
        RECT  0.16 2.24 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 2.80 0.28 ;
        RECT  2.34 -0.28 2.62 0.32 ;
        RECT  1.97 0.66 2.25 0.94 ;
        RECT  2.02 -0.28 2.18 0.94 ;
        END
    END GND!
END NAND4SP1V1_0

MACRO NAND4SP18V1_0
    CLASS CORE ;
    FOREIGN NAND4SP18V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.42 0.38 1.84 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.87 1.42 1.15 1.84 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.32 1.42 1.63 1.84 ;
        END
    END IN3
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.11 1.74 2.39 2.16 ;
        END
    END IN4
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 8.58  LAYER ME1  ;
        ANTENNADIFFAREA 5.25  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.58  LAYER ME1  ;
        ANTENNAMAXAREACAR 14.90  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.82 1.52 4.28 1.68 ;
        RECT  3.70 1.84 3.98 2.64 ;
        RECT  3.82 0.44 3.98 2.64 ;
        RECT  3.70 0.44 3.98 1.24 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.80 3.48 ;
        RECT  4.22 1.84 4.50 2.64 ;
        RECT  4.28 1.84 4.44 3.48 ;
        RECT  3.18 2.16 3.46 2.44 ;
        RECT  3.24 2.16 3.40 3.48 ;
        RECT  2.18 2.32 2.46 2.60 ;
        RECT  2.24 2.32 2.40 3.48 ;
        RECT  1.14 2.32 1.42 2.60 ;
        RECT  1.20 2.32 1.36 3.48 ;
        RECT  0.16 2.88 0.46 3.48 ;
        RECT  0.10 2.32 0.38 2.60 ;
        RECT  0.16 2.32 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.80 0.28 ;
        RECT  4.22 0.44 4.50 1.24 ;
        RECT  4.28 -0.28 4.44 1.24 ;
        RECT  3.18 0.64 3.46 0.92 ;
        RECT  3.24 -0.28 3.40 0.92 ;
        RECT  1.97 0.66 2.25 0.94 ;
        RECT  2.03 -0.28 2.19 0.94 ;
        RECT  0.18 -0.28 0.46 0.32 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.31 0.66 0.59 0.94 ;
        RECT  0.43 0.66 0.59 1.26 ;
        RECT  0.43 1.10 1.95 1.26 ;
        RECT  1.79 1.40 3.12 1.56 ;
        RECT  2.84 1.40 3.12 1.68 ;
        RECT  1.79 1.10 1.95 2.16 ;
        RECT  0.74 2.00 1.95 2.16 ;
        RECT  1.66 2.00 1.82 2.60 ;
        RECT  0.74 2.00 0.90 2.60 ;
        RECT  0.62 2.32 0.90 2.60 ;
        RECT  1.66 2.32 1.94 2.60 ;
        RECT  2.66 0.44 2.94 1.24 ;
        RECT  2.66 1.08 3.44 1.24 ;
        RECT  3.28 1.40 3.66 1.68 ;
        RECT  3.28 1.08 3.44 2.00 ;
        RECT  2.66 1.84 3.44 2.00 ;
        RECT  2.66 1.84 2.94 2.64 ;
    END
END NAND4SP18V1_0

MACRO NAND3SP8V1_0
    CLASS CORE ;
    FOREIGN NAND3SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 9.56  LAYER ME1  ;
        ANTENNADIFFAREA 7.67  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.82 1.97 5.10 2.25 ;
        RECT  0.62 2.00 5.10 2.16 ;
        RECT  3.78 1.97 4.06 2.25 ;
        RECT  2.70 1.97 2.98 2.25 ;
        RECT  1.66 1.97 1.94 2.25 ;
        RECT  1.08 0.76 1.42 1.04 ;
        RECT  0.22 1.20 1.24 1.36 ;
        RECT  1.08 0.76 1.24 1.36 ;
        RECT  0.62 1.97 1.08 2.16 ;
        RECT  0.92 1.20 1.08 2.16 ;
        RECT  0.62 1.97 0.90 2.25 ;
        RECT  0.22 0.76 0.38 1.36 ;
        RECT  0.10 0.76 0.38 1.04 ;
        END
    END OUT
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.58  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.40 1.39 1.68 1.81 ;
        RECT  1.32 1.52 1.68 1.68 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.58  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.96 1.39 3.24 1.81 ;
        RECT  2.92 1.52 3.24 1.68 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.46  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.57 1.39 4.85 1.81 ;
        RECT  4.52 1.52 4.85 1.68 ;
        END
    END IN3
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 5.20 3.48 ;
        RECT  4.74 2.88 5.02 3.48 ;
        RECT  4.30 2.32 4.58 2.60 ;
        RECT  4.36 2.32 4.52 3.48 ;
        RECT  3.22 2.48 3.50 2.76 ;
        RECT  3.28 2.48 3.44 3.48 ;
        RECT  2.18 2.48 2.46 2.76 ;
        RECT  2.24 2.48 2.40 3.48 ;
        RECT  1.14 2.48 1.42 2.76 ;
        RECT  1.20 2.48 1.36 3.48 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  0.16 2.48 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 5.20 0.28 ;
        RECT  4.82 0.76 5.10 1.04 ;
        RECT  4.74 -0.28 5.02 0.32 ;
        RECT  4.82 -0.28 4.98 1.04 ;
        RECT  3.90 0.48 4.98 0.64 ;
        RECT  3.78 0.76 4.06 1.04 ;
        RECT  3.90 0.48 4.06 1.04 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.74 0.44 1.82 0.60 ;
        RECT  1.66 0.44 1.82 1.04 ;
        RECT  0.74 0.44 0.90 1.04 ;
        RECT  0.62 0.76 0.90 1.04 ;
        RECT  1.66 0.76 2.00 1.04 ;
        RECT  2.64 0.76 2.98 1.04 ;
        RECT  1.84 0.76 2.00 1.36 ;
        RECT  2.64 0.76 2.80 1.36 ;
        RECT  1.84 1.20 2.80 1.36 ;
        RECT  2.30 0.44 3.38 0.60 ;
        RECT  3.22 0.44 3.38 1.04 ;
        RECT  2.30 0.44 2.46 1.04 ;
        RECT  2.18 0.76 2.46 1.04 ;
        RECT  3.22 0.76 3.56 1.04 ;
        RECT  4.25 0.80 4.58 1.08 ;
        RECT  3.40 0.76 3.56 1.36 ;
        RECT  4.25 0.80 4.41 1.36 ;
        RECT  3.40 1.20 4.41 1.36 ;
    END
END NAND3SP8V1_0

MACRO NAND3SP5V1_0
    CLASS CORE ;
    FOREIGN NAND3SP5V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.38  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.40 0.58 1.68 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.38  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.46 1.32 2.74 1.74 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.34  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.49 1.46 3.91 1.74 ;
        END
    END IN3
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 7.96  LAYER ME1  ;
        ANTENNADIFFAREA 6.06  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.24 2.22 3.52 2.50 ;
        RECT  3.24 1.92 3.40 2.50 ;
        RECT  0.76 1.92 3.40 2.08 ;
        RECT  1.68 2.24 1.96 2.52 ;
        RECT  1.74 1.92 1.90 2.52 ;
        RECT  0.64 2.22 0.92 2.50 ;
        RECT  0.76 0.76 0.92 2.50 ;
        RECT  0.64 0.76 0.92 1.04 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.40 3.48 ;
        RECT  3.82 2.88 4.22 3.48 ;
        RECT  3.76 2.38 4.04 2.66 ;
        RECT  3.82 2.38 3.98 3.48 ;
        RECT  2.72 2.38 3.00 2.66 ;
        RECT  2.78 2.38 2.94 3.48 ;
        RECT  2.20 2.48 2.48 2.76 ;
        RECT  2.26 2.48 2.42 3.48 ;
        RECT  1.16 2.48 1.44 2.76 ;
        RECT  1.22 2.48 1.38 3.48 ;
        RECT  0.12 2.48 0.40 2.76 ;
        RECT  0.18 2.48 0.34 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.40 0.28 ;
        RECT  3.94 -0.28 4.22 0.32 ;
        RECT  3.24 0.70 3.52 0.98 ;
        RECT  3.26 -0.28 3.42 0.98 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.24 0.44 1.32 0.60 ;
        RECT  0.24 0.44 0.40 1.04 ;
        RECT  0.12 0.76 0.40 1.04 ;
        RECT  1.16 0.44 1.32 1.04 ;
        RECT  2.14 0.76 2.48 1.04 ;
        RECT  1.28 0.76 1.44 1.36 ;
        RECT  2.14 0.76 2.30 1.36 ;
        RECT  1.28 1.20 2.30 1.36 ;
        RECT  1.80 0.44 2.88 0.60 ;
        RECT  2.72 0.44 2.88 0.98 ;
        RECT  2.72 0.70 3.06 0.98 ;
        RECT  3.76 0.70 4.04 0.98 ;
        RECT  1.80 0.44 1.96 1.04 ;
        RECT  1.68 0.76 1.96 1.04 ;
        RECT  2.90 0.70 3.06 1.30 ;
        RECT  3.76 0.70 3.92 1.30 ;
        RECT  2.90 1.14 3.92 1.30 ;
    END
END NAND3SP5V1_0

MACRO NAND3SP2V1_0
    CLASS CORE ;
    FOREIGN NAND3SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 2.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.14  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.14  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.34 1.14 1.76 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.14  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.34 1.34 1.62 1.76 ;
        RECT  1.32 1.52 1.62 1.68 ;
        END
    END IN3
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 3.07  LAYER ME1  ;
        ANTENNADIFFAREA 2.51  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.66 2.06 1.94 2.34 ;
        RECT  0.54 1.92 1.82 2.08 ;
        RECT  0.62 1.92 0.90 2.34 ;
        RECT  0.54 0.96 0.70 2.08 ;
        RECT  0.24 0.96 0.70 1.12 ;
        RECT  0.24 0.84 0.52 1.12 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 2.40 3.48 ;
        RECT  1.94 2.88 2.22 3.48 ;
        RECT  1.14 2.38 1.42 2.66 ;
        RECT  1.20 2.38 1.36 3.48 ;
        RECT  0.10 2.38 0.38 2.66 ;
        RECT  0.16 2.38 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 2.40 0.28 ;
        RECT  1.94 -0.28 2.22 0.32 ;
        RECT  1.52 0.52 1.80 0.80 ;
        RECT  1.58 -0.28 1.74 0.80 ;
        END
    END GND!
END NAND3SP2V1_0

MACRO NAND3SP1V1_0
    CLASS CORE ;
    FOREIGN NAND3SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 2.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.44 1.32 0.72 1.74 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.92 1.32 1.20 1.74 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.48 1.46 1.94 1.74 ;
        END
    END IN3
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 3.17  LAYER ME1  ;
        ANTENNADIFFAREA 1.76  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.14 2.22 1.42 2.50 ;
        RECT  1.16 1.90 1.32 2.50 ;
        RECT  0.12 1.90 1.32 2.06 ;
        RECT  0.12 0.80 0.50 1.08 ;
        RECT  0.10 2.22 0.38 2.50 ;
        RECT  0.12 0.80 0.28 2.50 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 2.40 3.48 ;
        RECT  1.72 2.88 2.22 3.48 ;
        RECT  1.66 2.22 1.94 2.50 ;
        RECT  1.72 2.22 1.88 3.48 ;
        RECT  0.62 2.22 0.90 2.50 ;
        RECT  0.68 2.22 0.84 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 2.40 0.28 ;
        RECT  1.94 -0.28 2.22 0.32 ;
        RECT  1.50 0.80 1.78 1.08 ;
        RECT  1.54 -0.28 1.70 1.08 ;
        END
    END GND!
END NAND3SP1V1_0

MACRO NAND3SP14V1_0
    CLASS CORE ;
    FOREIGN NAND3SP14V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.96  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.39 1.46 2.77 1.74 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.96  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.86 1.46 5.32 1.74 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.96  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.66 1.32 7.94 1.74 ;
        END
    END IN3
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 16.78  LAYER ME1  ;
        ANTENNADIFFAREA 13.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.90 2.22 8.18 2.50 ;
        RECT  7.94 1.90 8.10 2.50 ;
        RECT  0.74 1.90 8.10 2.06 ;
        RECT  6.86 2.22 7.14 2.50 ;
        RECT  6.92 1.90 7.08 2.50 ;
        RECT  5.82 2.22 6.10 2.50 ;
        RECT  5.88 1.90 6.04 2.50 ;
        RECT  4.78 2.22 5.06 2.50 ;
        RECT  4.84 1.90 5.00 2.50 ;
        RECT  3.74 2.22 4.02 2.50 ;
        RECT  3.80 1.90 3.96 2.50 ;
        RECT  2.70 2.22 2.98 2.50 ;
        RECT  2.76 1.90 2.92 2.50 ;
        RECT  2.10 0.76 2.46 1.04 ;
        RECT  0.22 1.20 2.26 1.36 ;
        RECT  2.10 0.76 2.26 1.36 ;
        RECT  1.66 2.22 1.94 2.50 ;
        RECT  1.72 1.90 1.88 2.50 ;
        RECT  1.32 1.20 1.48 2.06 ;
        RECT  1.14 0.76 1.42 1.04 ;
        RECT  1.20 0.76 1.36 1.36 ;
        RECT  0.62 2.22 0.90 2.50 ;
        RECT  0.74 1.90 0.90 2.50 ;
        RECT  0.22 0.76 0.38 1.36 ;
        RECT  0.10 0.76 0.38 1.04 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 9.20 3.48 ;
        RECT  8.74 2.88 9.02 3.48 ;
        RECT  7.38 2.48 7.66 2.76 ;
        RECT  7.44 2.48 7.60 3.48 ;
        RECT  6.34 2.48 6.62 2.76 ;
        RECT  6.40 2.48 6.56 3.48 ;
        RECT  5.30 2.48 5.58 2.76 ;
        RECT  5.36 2.48 5.52 3.48 ;
        RECT  4.26 2.48 4.54 2.76 ;
        RECT  4.32 2.48 4.48 3.48 ;
        RECT  3.22 2.48 3.50 2.76 ;
        RECT  3.28 2.48 3.44 3.48 ;
        RECT  2.18 2.48 2.46 2.76 ;
        RECT  2.24 2.48 2.40 3.48 ;
        RECT  1.14 2.48 1.42 2.76 ;
        RECT  1.20 2.48 1.36 3.48 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  0.16 2.48 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 9.20 0.28 ;
        RECT  8.74 -0.28 9.02 0.32 ;
        RECT  7.90 0.76 8.18 1.04 ;
        RECT  7.96 -0.28 8.12 1.04 ;
        RECT  6.86 0.76 7.14 1.04 ;
        RECT  6.92 -0.28 7.08 1.04 ;
        RECT  5.82 0.76 6.10 1.04 ;
        RECT  5.88 -0.28 6.04 1.04 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.74 0.44 2.86 0.60 ;
        RECT  1.72 0.44 1.88 1.04 ;
        RECT  2.70 0.44 2.86 1.04 ;
        RECT  0.74 0.44 0.90 1.04 ;
        RECT  0.62 0.76 0.90 1.04 ;
        RECT  1.66 0.76 1.94 1.04 ;
        RECT  2.70 0.76 3.06 1.04 ;
        RECT  3.74 0.76 4.02 1.04 ;
        RECT  4.78 0.76 5.06 1.04 ;
        RECT  4.47 0.88 5.06 1.04 ;
        RECT  2.90 0.76 3.06 1.36 ;
        RECT  3.80 0.76 3.96 1.36 ;
        RECT  4.47 0.88 4.63 1.36 ;
        RECT  2.90 1.20 4.63 1.36 ;
        RECT  3.34 0.44 5.46 0.60 ;
        RECT  4.26 0.44 4.54 0.72 ;
        RECT  5.30 0.44 5.46 1.04 ;
        RECT  3.34 0.44 3.50 1.04 ;
        RECT  3.22 0.76 3.50 1.04 ;
        RECT  5.30 0.76 5.64 1.04 ;
        RECT  6.34 0.76 6.62 1.04 ;
        RECT  7.32 0.76 7.66 1.04 ;
        RECT  5.48 0.76 5.64 1.36 ;
        RECT  6.40 0.76 6.56 1.36 ;
        RECT  7.32 0.76 7.48 1.36 ;
        RECT  5.48 1.20 7.48 1.36 ;
    END
END NAND3SP14V1_0

MACRO NAND2SP9V1_0
    CLASS CORE ;
    FOREIGN NAND2SP9V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.43  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.26 1.52 0.68 1.80 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.43  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.86 1.47 3.28 1.75 ;
        END
    END IN2
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 6.74  LAYER ME1  ;
        ANTENNADIFFAREA 4.74  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.70 2.21 2.98 2.49 ;
        RECT  2.70 1.91 2.86 2.49 ;
        RECT  0.80 1.91 2.86 2.07 ;
        RECT  1.66 2.23 1.94 2.51 ;
        RECT  1.72 1.91 1.88 2.51 ;
        RECT  1.20 1.52 1.48 1.68 ;
        RECT  1.14 0.76 1.42 1.04 ;
        RECT  1.20 0.76 1.36 2.07 ;
        RECT  0.22 1.20 1.36 1.36 ;
        RECT  0.62 2.21 0.96 2.49 ;
        RECT  0.80 1.91 0.96 2.49 ;
        RECT  0.22 0.76 0.38 1.36 ;
        RECT  0.10 0.76 0.38 1.04 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 3.60 3.48 ;
        RECT  3.22 2.21 3.50 2.49 ;
        RECT  3.14 2.88 3.44 3.48 ;
        RECT  3.28 2.21 3.44 3.48 ;
        RECT  2.18 2.23 2.46 2.51 ;
        RECT  2.24 2.23 2.40 3.48 ;
        RECT  1.14 2.23 1.42 2.51 ;
        RECT  1.20 2.23 1.36 3.48 ;
        RECT  0.10 2.21 0.38 2.49 ;
        RECT  0.16 2.21 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 3.60 0.28 ;
        RECT  3.22 0.71 3.50 0.99 ;
        RECT  3.28 -0.28 3.44 0.99 ;
        RECT  3.14 -0.28 3.44 0.32 ;
        RECT  2.18 0.71 2.46 0.99 ;
        RECT  2.24 -0.28 2.40 0.99 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.74 0.44 1.82 0.60 ;
        RECT  2.70 0.71 2.98 0.99 ;
        RECT  0.74 0.44 0.90 1.04 ;
        RECT  0.62 0.76 0.90 1.04 ;
        RECT  1.66 0.44 1.82 1.04 ;
        RECT  1.78 0.76 1.94 1.31 ;
        RECT  2.70 0.71 2.86 1.31 ;
        RECT  1.78 1.15 2.86 1.31 ;
    END
END NAND2SP9V1_0

MACRO NAND2SP6V1_0
    CLASS CORE ;
    FOREIGN NAND2SP6V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 2.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.29  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.32 1.46 0.74 1.74 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.29  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.12 1.52 2.54 1.81 ;
        END
    END IN2
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 4.51  LAYER ME1  ;
        ANTENNADIFFAREA 3.57  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.80 2.07 2.10 2.36 ;
        RECT  1.80 1.75 1.96 2.36 ;
        RECT  0.92 1.75 1.96 1.91 ;
        RECT  0.78 2.07 1.08 2.36 ;
        RECT  0.92 0.76 1.08 2.36 ;
        RECT  0.78 0.76 1.08 1.05 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 2.80 3.48 ;
        RECT  2.34 2.88 2.62 3.48 ;
        RECT  2.34 2.07 2.62 2.36 ;
        RECT  2.40 2.07 2.56 3.48 ;
        RECT  1.30 2.07 1.58 2.36 ;
        RECT  1.36 2.07 1.52 3.48 ;
        RECT  0.26 2.07 0.54 2.36 ;
        RECT  0.32 2.07 0.48 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 2.80 0.28 ;
        RECT  2.34 -0.28 2.62 0.32 ;
        RECT  1.82 0.75 2.10 1.04 ;
        RECT  1.88 -0.28 2.04 1.04 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.38 0.44 1.46 0.60 ;
        RECT  1.30 0.44 1.46 1.04 ;
        RECT  2.34 0.75 2.62 1.04 ;
        RECT  0.38 0.44 0.54 1.05 ;
        RECT  0.26 0.76 0.54 1.05 ;
        RECT  1.42 0.75 1.58 1.36 ;
        RECT  2.34 0.75 2.50 1.36 ;
        RECT  1.42 1.20 2.50 1.36 ;
    END
END NAND2SP6V1_0

MACRO NAND2SP3V1_0
    CLASS CORE ;
    FOREIGN NAND2SP3V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 1.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.15  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.46 0.52 1.74 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.15  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.00 1.46 1.52 1.74 ;
        END
    END IN2
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 2.49  LAYER ME1  ;
        ANTENNADIFFAREA 1.90  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.62 1.94 0.90 2.56 ;
        RECT  0.68 1.08 0.84 2.56 ;
        RECT  0.49 1.08 0.84 1.28 ;
        RECT  0.17 1.08 0.84 1.24 ;
        RECT  0.17 0.62 0.45 1.24 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 1.60 3.48 ;
        RECT  1.14 2.88 1.42 3.48 ;
        RECT  1.14 1.94 1.42 2.56 ;
        RECT  1.20 1.94 1.36 3.48 ;
        RECT  0.10 1.94 0.38 2.56 ;
        RECT  0.16 1.94 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 1.60 0.28 ;
        RECT  1.13 -0.28 1.42 0.32 ;
        RECT  1.07 0.62 1.35 1.24 ;
        RECT  1.13 -0.28 1.29 1.24 ;
        END
    END GND!
END NAND2SP3V1_0

MACRO NAND2SP2V1_0
    CLASS CORE ;
    FOREIGN NAND2SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 1.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 2.32  LAYER ME1  ;
        ANTENNADIFFAREA 1.45  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.54 1.92 0.90 2.20 ;
        RECT  0.54 1.08 0.70 2.20 ;
        RECT  0.52 1.08 0.70 1.28 ;
        RECT  0.10 1.08 0.70 1.24 ;
        RECT  0.10 0.96 0.38 1.24 ;
        END
    END OUT
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.10  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.46 0.38 1.88 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.10  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.34 1.14 1.76 ;
        END
    END IN2
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 1.60 3.48 ;
        RECT  1.14 2.88 1.42 3.48 ;
        RECT  1.14 2.04 1.42 2.32 ;
        RECT  1.20 2.04 1.36 3.48 ;
        RECT  0.10 2.04 0.38 2.32 ;
        RECT  0.16 2.04 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 1.60 0.28 ;
        RECT  1.06 -0.28 1.42 0.32 ;
        RECT  1.00 0.84 1.28 1.12 ;
        RECT  1.06 -0.28 1.22 1.12 ;
        END
    END GND!
END NAND2SP2V1_0

MACRO NAND2SP28V1_0
    CLASS CORE ;
    FOREIGN NAND2SP28V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.31  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.32 1.46 0.74 1.74 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.31  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.38 1.46 8.80 1.74 ;
        END
    END IN2
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 17.72  LAYER ME1  ;
        ANTENNADIFFAREA 12.44  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.06 2.09 8.34 2.37 ;
        RECT  8.06 1.77 8.22 2.37 ;
        RECT  0.90 1.77 8.22 1.93 ;
        RECT  7.02 2.09 7.30 2.37 ;
        RECT  7.08 1.77 7.24 2.37 ;
        RECT  5.98 2.09 6.26 2.37 ;
        RECT  6.04 1.77 6.20 2.37 ;
        RECT  4.94 2.09 5.22 2.37 ;
        RECT  5.00 1.77 5.16 2.37 ;
        RECT  3.90 2.09 4.18 2.37 ;
        RECT  3.90 0.76 4.18 1.04 ;
        RECT  3.96 1.77 4.12 2.37 ;
        RECT  0.90 1.20 4.06 1.36 ;
        RECT  3.90 0.76 4.06 1.36 ;
        RECT  2.86 2.09 3.14 2.37 ;
        RECT  2.86 0.76 3.14 1.04 ;
        RECT  2.92 1.77 3.08 2.37 ;
        RECT  2.92 0.76 3.08 1.36 ;
        RECT  2.52 1.20 2.68 1.93 ;
        RECT  1.82 2.09 2.10 2.37 ;
        RECT  1.82 0.76 2.10 1.04 ;
        RECT  1.88 1.77 2.04 2.37 ;
        RECT  1.88 0.76 2.04 1.36 ;
        RECT  0.78 2.09 1.06 2.37 ;
        RECT  0.90 1.77 1.06 2.37 ;
        RECT  0.90 0.76 1.06 1.36 ;
        RECT  0.78 0.76 1.06 1.04 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 9.20 3.48 ;
        RECT  8.64 2.88 9.02 3.48 ;
        RECT  8.58 2.09 8.86 2.37 ;
        RECT  8.64 2.09 8.80 3.48 ;
        RECT  7.54 2.09 7.82 2.37 ;
        RECT  7.60 2.09 7.76 3.48 ;
        RECT  6.50 2.09 6.78 2.37 ;
        RECT  6.56 2.09 6.72 3.48 ;
        RECT  5.46 2.09 5.74 2.37 ;
        RECT  5.52 2.09 5.68 3.48 ;
        RECT  4.42 2.09 4.70 2.37 ;
        RECT  4.48 2.09 4.64 3.48 ;
        RECT  3.38 2.09 3.66 2.37 ;
        RECT  3.44 2.09 3.60 3.48 ;
        RECT  2.34 2.09 2.62 2.37 ;
        RECT  2.40 2.09 2.56 3.48 ;
        RECT  1.30 2.09 1.58 2.37 ;
        RECT  1.36 2.09 1.52 3.48 ;
        RECT  0.26 2.09 0.54 2.37 ;
        RECT  0.32 2.09 0.48 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 9.20 0.28 ;
        RECT  8.74 -0.28 9.02 0.32 ;
        RECT  8.06 0.70 8.34 0.98 ;
        RECT  8.12 -0.28 8.28 0.98 ;
        RECT  7.02 0.75 7.30 1.03 ;
        RECT  7.08 -0.28 7.24 1.03 ;
        RECT  5.98 0.75 6.26 1.03 ;
        RECT  6.04 -0.28 6.20 1.03 ;
        RECT  4.94 0.75 5.22 1.03 ;
        RECT  5.00 -0.28 5.16 1.03 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.38 0.44 4.58 0.60 ;
        RECT  1.36 0.44 1.52 1.04 ;
        RECT  2.40 0.44 2.56 1.04 ;
        RECT  3.44 0.44 3.60 1.04 ;
        RECT  7.54 0.70 7.82 0.98 ;
        RECT  4.42 0.44 4.58 1.03 ;
        RECT  5.46 0.75 5.74 1.03 ;
        RECT  6.50 0.75 6.78 1.03 ;
        RECT  0.38 0.44 0.54 1.04 ;
        RECT  0.26 0.76 0.54 1.04 ;
        RECT  1.30 0.76 1.58 1.04 ;
        RECT  2.34 0.76 2.62 1.04 ;
        RECT  3.38 0.76 3.66 1.04 ;
        RECT  8.58 0.76 8.86 1.04 ;
        RECT  4.54 0.75 4.70 1.35 ;
        RECT  5.52 0.75 5.68 1.35 ;
        RECT  6.56 0.75 6.72 1.35 ;
        RECT  7.60 1.14 8.74 1.30 ;
        RECT  8.58 0.76 8.74 1.30 ;
        RECT  7.60 0.70 7.76 1.35 ;
        RECT  4.54 1.19 7.76 1.35 ;
    END
END NAND2SP28V1_0

MACRO NAND2SP1V1_0
    CLASS CORE ;
    FOREIGN NAND2SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 1.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.40 0.38 1.82 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.40 1.14 1.82 ;
        END
    END IN2
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 2.36  LAYER ME1  ;
        ANTENNADIFFAREA 1.21  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.54 1.98 0.90 2.26 ;
        RECT  0.54 1.08 0.70 2.26 ;
        RECT  0.52 1.08 0.70 1.28 ;
        RECT  0.10 1.08 0.70 1.24 ;
        RECT  0.10 0.96 0.38 1.24 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 1.60 3.48 ;
        RECT  1.14 2.88 1.42 3.48 ;
        RECT  1.14 1.98 1.42 2.26 ;
        RECT  1.20 1.98 1.36 3.48 ;
        RECT  0.10 1.98 0.38 2.26 ;
        RECT  0.16 1.98 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 1.60 0.28 ;
        RECT  1.06 -0.28 1.42 0.32 ;
        RECT  1.00 0.96 1.28 1.24 ;
        RECT  1.06 -0.28 1.22 1.24 ;
        END
    END GND!
END NAND2SP1V1_0

MACRO NAND2SP14V1_0
    CLASS CORE ;
    FOREIGN NAND2SP14V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.26 1.40 0.68 1.68 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.06 1.46 4.48 1.74 ;
        END
    END IN2
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 9.00  LAYER ME1  ;
        ANTENNADIFFAREA 6.82  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.78 2.16 4.06 2.44 ;
        RECT  3.78 1.88 3.94 2.44 ;
        RECT  2.86 1.88 3.94 2.04 ;
        RECT  2.74 2.16 3.02 2.44 ;
        RECT  2.86 1.83 3.02 2.44 ;
        RECT  0.78 1.83 3.02 1.99 ;
        RECT  1.70 2.16 1.98 2.44 ;
        RECT  1.70 0.76 1.98 1.04 ;
        RECT  1.76 1.83 1.92 2.44 ;
        RECT  0.78 1.11 1.86 1.27 ;
        RECT  1.70 0.76 1.86 1.27 ;
        RECT  1.32 1.11 1.48 1.99 ;
        RECT  0.66 2.16 0.94 2.44 ;
        RECT  0.78 1.83 0.94 2.44 ;
        RECT  0.78 0.76 0.94 1.27 ;
        RECT  0.66 0.76 0.94 1.04 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.80 3.48 ;
        RECT  4.34 2.88 4.62 3.48 ;
        RECT  4.30 2.16 4.58 2.44 ;
        RECT  4.36 2.16 4.52 3.48 ;
        RECT  3.26 2.21 3.54 2.49 ;
        RECT  3.32 2.21 3.48 3.48 ;
        RECT  2.22 2.16 2.50 2.44 ;
        RECT  2.28 2.16 2.44 3.48 ;
        RECT  1.18 2.16 1.46 2.44 ;
        RECT  1.24 2.16 1.40 3.48 ;
        RECT  0.14 2.16 0.42 2.44 ;
        RECT  0.20 2.16 0.36 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.80 0.28 ;
        RECT  4.34 -0.28 4.62 0.32 ;
        RECT  3.78 0.66 4.06 0.94 ;
        RECT  3.88 -0.28 4.04 0.94 ;
        RECT  2.74 0.71 3.02 0.99 ;
        RECT  2.84 -0.28 3.00 0.99 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.26 0.44 2.38 0.60 ;
        RECT  1.18 0.44 1.46 0.95 ;
        RECT  2.22 0.44 2.38 0.99 ;
        RECT  3.26 0.71 3.54 0.99 ;
        RECT  4.30 0.71 4.58 0.99 ;
        RECT  0.26 0.44 0.42 1.00 ;
        RECT  0.14 0.72 0.42 1.00 ;
        RECT  2.34 0.71 2.50 1.31 ;
        RECT  3.38 1.10 4.46 1.26 ;
        RECT  4.30 0.71 4.46 1.26 ;
        RECT  3.38 0.71 3.54 1.31 ;
        RECT  2.34 1.15 3.54 1.31 ;
    END
END NAND2SP14V1_0

MACRO MUX5SP8V1_0
    CLASS CORE ;
    FOREIGN MUX5SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 24.34  LAYER ME1  ;
        ANTENNADIFFAREA 11.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.11  LAYER ME1  ;
        ANTENNAMAXAREACAR 21.95  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.64 1.84 13.92 2.12 ;
        RECT  13.64 0.96 13.92 1.24 ;
        RECT  13.64 0.96 13.80 2.12 ;
        RECT  11.72 1.52 13.80 1.68 ;
        RECT  12.60 1.84 12.88 2.12 ;
        RECT  12.60 0.96 12.88 1.24 ;
        RECT  12.66 0.96 12.82 2.12 ;
        RECT  11.56 1.84 11.88 2.12 ;
        RECT  11.72 0.96 11.88 2.12 ;
        RECT  11.56 0.96 11.88 1.24 ;
        END
    END OUT
    PIN S2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.68 1.38 11.08 1.68 ;
        END
    END S2
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.60 1.26 7.88 1.68 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.46 0.50 1.74 ;
        END
    END S0
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.08 1.26 8.36 1.68 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.33  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 19.73  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.66 0.76 3.94 2.20 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.96  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 14.21  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.76 1.46 3.14 1.74 ;
        RECT  2.62 1.92 2.92 2.20 ;
        RECT  2.76 0.76 2.92 2.20 ;
        RECT  2.62 0.76 2.92 1.04 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.49  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 22.12  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.14 1.92 2.42 2.20 ;
        RECT  2.14 0.76 2.42 1.04 ;
        RECT  2.14 0.76 2.34 2.20 ;
        RECT  2.06 1.46 2.34 1.74 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.14  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.02  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.22 1.46 1.54 1.74 ;
        RECT  1.10 1.92 1.38 2.20 ;
        RECT  1.22 0.76 1.38 2.20 ;
        RECT  1.10 0.76 1.38 1.04 ;
        END
    END A
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 14.40 3.48 ;
        RECT  13.94 2.88 14.22 3.48 ;
        RECT  13.12 2.26 13.40 2.54 ;
        RECT  13.18 2.26 13.34 3.48 ;
        RECT  12.08 2.26 12.36 2.54 ;
        RECT  12.14 2.26 12.30 3.48 ;
        RECT  10.95 2.62 11.23 3.48 ;
        RECT  7.82 2.62 8.10 3.48 ;
        RECT  4.59 2.62 4.87 3.48 ;
        RECT  0.10 1.90 0.38 2.18 ;
        RECT  0.16 1.90 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 14.40 0.28 ;
        RECT  13.94 -0.28 14.22 0.32 ;
        RECT  13.12 0.54 13.40 0.82 ;
        RECT  13.18 -0.28 13.34 0.82 ;
        RECT  12.08 0.54 12.36 0.82 ;
        RECT  12.14 -0.28 12.30 0.82 ;
        RECT  11.04 0.94 11.32 1.22 ;
        RECT  11.10 -0.28 11.26 1.22 ;
        RECT  7.78 0.82 8.06 1.10 ;
        RECT  7.84 -0.28 8.00 1.10 ;
        RECT  4.76 0.96 5.04 1.24 ;
        RECT  4.82 -0.28 4.98 1.24 ;
        RECT  0.10 0.96 0.38 1.24 ;
        RECT  0.16 -0.28 0.32 1.24 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.96 0.90 1.24 ;
        RECT  0.68 1.40 1.04 1.68 ;
        RECT  0.68 0.96 0.84 2.18 ;
        RECT  0.62 1.90 0.90 2.18 ;
        RECT  3.30 0.44 4.38 0.60 ;
        RECT  4.10 0.44 4.38 0.72 ;
        RECT  3.14 0.76 3.46 1.04 ;
        RECT  3.30 0.44 3.46 2.20 ;
        RECT  3.14 1.92 3.46 2.20 ;
        RECT  1.62 0.76 1.90 1.04 ;
        RECT  1.70 0.76 1.86 2.20 ;
        RECT  1.62 1.92 1.90 2.20 ;
        RECT  1.74 1.92 1.90 2.52 ;
        RECT  1.74 2.36 4.44 2.52 ;
        RECT  4.16 2.28 4.44 2.56 ;
        RECT  5.32 0.76 5.60 1.04 ;
        RECT  5.38 0.76 5.54 2.20 ;
        RECT  5.32 1.92 5.60 2.20 ;
        RECT  6.34 0.76 6.64 1.04 ;
        RECT  4.24 0.96 4.52 1.24 ;
        RECT  4.30 0.96 4.46 2.12 ;
        RECT  6.34 0.76 6.50 2.20 ;
        RECT  4.24 1.84 4.52 2.12 ;
        RECT  4.24 1.96 5.16 2.12 ;
        RECT  6.34 1.92 6.64 2.20 ;
        RECT  5.00 1.96 5.16 2.52 ;
        RECT  6.36 1.92 6.52 2.52 ;
        RECT  5.00 2.36 6.52 2.52 ;
        RECT  7.26 0.82 7.54 1.10 ;
        RECT  7.12 1.40 7.42 1.68 ;
        RECT  7.26 0.82 7.42 2.12 ;
        RECT  7.26 1.84 7.54 2.12 ;
        RECT  5.96 0.44 6.96 0.60 ;
        RECT  5.96 0.44 6.12 1.04 ;
        RECT  5.84 0.76 6.12 1.04 ;
        RECT  8.88 0.76 9.16 1.04 ;
        RECT  5.90 0.76 6.06 2.20 ;
        RECT  8.94 0.76 9.10 2.20 ;
        RECT  5.84 1.92 6.12 2.20 ;
        RECT  8.88 1.92 9.16 2.20 ;
        RECT  6.80 0.44 6.96 2.44 ;
        RECT  8.88 1.92 9.04 2.44 ;
        RECT  6.80 2.28 9.04 2.44 ;
        RECT  8.52 0.44 10.08 0.60 ;
        RECT  9.92 0.76 10.20 1.04 ;
        RECT  8.30 0.82 8.68 1.10 ;
        RECT  9.92 0.44 10.08 2.20 ;
        RECT  8.52 0.44 8.68 2.12 ;
        RECT  8.30 1.84 8.68 2.12 ;
        RECT  9.92 1.92 10.20 2.20 ;
        RECT  10.36 0.94 10.80 1.22 ;
        RECT  10.24 1.40 10.52 1.68 ;
        RECT  10.36 0.94 10.52 2.12 ;
        RECT  10.36 1.84 10.80 2.12 ;
        RECT  9.40 0.76 9.68 1.04 ;
        RECT  11.24 1.40 11.56 1.68 ;
        RECT  9.46 0.76 9.62 2.20 ;
        RECT  9.40 1.92 9.68 2.20 ;
        RECT  9.52 1.92 9.68 2.52 ;
        RECT  10.52 2.28 11.40 2.44 ;
        RECT  11.24 1.40 11.40 2.44 ;
        RECT  9.52 2.36 10.68 2.52 ;
    END
END MUX5SP8V1_0

MACRO MUX5SP4V1_0
    CLASS CORE ;
    FOREIGN MUX5SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.14  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.02  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.22 1.46 1.54 1.74 ;
        RECT  1.10 1.92 1.38 2.20 ;
        RECT  1.22 0.76 1.38 2.20 ;
        RECT  1.10 0.76 1.38 1.04 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.49  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 22.12  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.14 1.92 2.42 2.20 ;
        RECT  2.14 0.76 2.42 1.04 ;
        RECT  2.14 0.76 2.34 2.20 ;
        RECT  2.06 1.46 2.34 1.74 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.96  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 14.21  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.76 1.46 3.14 1.74 ;
        RECT  2.62 1.92 2.92 2.20 ;
        RECT  2.76 0.76 2.92 2.20 ;
        RECT  2.62 0.76 2.92 1.04 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.33  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 19.73  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.66 0.76 3.94 2.20 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.08 1.26 8.36 1.68 ;
        END
    END E
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.46 0.50 1.74 ;
        END
    END S0
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.60 1.26 7.88 1.68 ;
        END
    END S1
    PIN S2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.68 1.38 11.08 1.68 ;
        END
    END S2
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 21.28  LAYER ME1  ;
        ANTENNADIFFAREA 9.26  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER ME1  ;
        ANTENNAMAXAREACAR 37.57  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.56 1.84 11.88 2.12 ;
        RECT  11.72 0.94 11.88 2.12 ;
        RECT  11.56 0.94 11.88 1.22 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 12.80 3.48 ;
        RECT  12.14 2.88 12.62 3.48 ;
        RECT  12.08 2.18 12.36 2.46 ;
        RECT  12.14 2.18 12.30 3.48 ;
        RECT  10.95 2.62 11.23 3.48 ;
        RECT  7.82 2.62 8.10 3.48 ;
        RECT  4.59 2.62 4.87 3.48 ;
        RECT  0.10 1.90 0.38 2.18 ;
        RECT  0.16 1.90 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 12.80 0.28 ;
        RECT  12.14 -0.28 12.62 0.32 ;
        RECT  12.08 0.60 12.36 0.88 ;
        RECT  12.14 -0.28 12.30 0.88 ;
        RECT  11.04 0.94 11.32 1.22 ;
        RECT  11.10 -0.28 11.26 1.22 ;
        RECT  7.78 0.82 8.06 1.10 ;
        RECT  7.84 -0.28 8.00 1.10 ;
        RECT  4.76 0.96 5.04 1.24 ;
        RECT  4.82 -0.28 4.98 1.24 ;
        RECT  0.10 0.96 0.38 1.24 ;
        RECT  0.16 -0.28 0.32 1.24 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.96 0.90 1.24 ;
        RECT  0.68 1.40 1.04 1.68 ;
        RECT  0.68 0.96 0.84 2.18 ;
        RECT  0.62 1.90 0.90 2.18 ;
        RECT  3.30 0.44 4.38 0.60 ;
        RECT  4.10 0.44 4.38 0.72 ;
        RECT  3.14 0.76 3.46 1.04 ;
        RECT  3.30 0.44 3.46 2.20 ;
        RECT  3.14 1.92 3.46 2.20 ;
        RECT  1.62 0.76 1.90 1.04 ;
        RECT  1.70 0.76 1.86 2.20 ;
        RECT  1.62 1.92 1.90 2.20 ;
        RECT  1.74 1.92 1.90 2.52 ;
        RECT  1.74 2.36 4.44 2.52 ;
        RECT  4.16 2.28 4.44 2.56 ;
        RECT  5.32 0.76 5.60 1.04 ;
        RECT  5.38 0.76 5.54 2.20 ;
        RECT  5.32 1.92 5.60 2.20 ;
        RECT  6.34 0.76 6.64 1.04 ;
        RECT  4.24 0.96 4.52 1.24 ;
        RECT  4.30 0.96 4.46 2.12 ;
        RECT  6.34 0.76 6.50 2.20 ;
        RECT  4.24 1.84 4.52 2.12 ;
        RECT  4.24 1.96 5.16 2.12 ;
        RECT  6.34 1.92 6.64 2.20 ;
        RECT  5.00 1.96 5.16 2.52 ;
        RECT  6.36 1.92 6.52 2.52 ;
        RECT  5.00 2.36 6.52 2.52 ;
        RECT  7.26 0.82 7.54 1.10 ;
        RECT  7.12 1.40 7.42 1.68 ;
        RECT  7.26 0.82 7.42 2.12 ;
        RECT  7.26 1.84 7.54 2.12 ;
        RECT  5.96 0.44 6.96 0.60 ;
        RECT  5.96 0.44 6.12 1.04 ;
        RECT  5.84 0.76 6.12 1.04 ;
        RECT  8.88 0.76 9.16 1.04 ;
        RECT  5.90 0.76 6.06 2.20 ;
        RECT  8.94 0.76 9.10 2.20 ;
        RECT  5.84 1.92 6.12 2.20 ;
        RECT  8.88 1.92 9.16 2.20 ;
        RECT  6.80 0.44 6.96 2.44 ;
        RECT  8.88 1.92 9.04 2.44 ;
        RECT  6.80 2.28 9.04 2.44 ;
        RECT  8.52 0.44 10.08 0.60 ;
        RECT  9.92 0.76 10.20 1.04 ;
        RECT  8.30 0.82 8.68 1.10 ;
        RECT  9.92 0.44 10.08 2.20 ;
        RECT  8.52 0.44 8.68 2.12 ;
        RECT  8.30 1.84 8.68 2.12 ;
        RECT  9.92 1.92 10.20 2.20 ;
        RECT  10.36 0.94 10.80 1.22 ;
        RECT  10.24 1.40 10.52 1.68 ;
        RECT  10.36 0.94 10.52 2.12 ;
        RECT  10.36 1.84 10.80 2.12 ;
        RECT  9.40 0.76 9.68 1.04 ;
        RECT  11.24 1.40 11.56 1.68 ;
        RECT  9.46 0.76 9.62 2.20 ;
        RECT  9.40 1.92 9.68 2.20 ;
        RECT  9.52 1.92 9.68 2.52 ;
        RECT  10.52 2.28 11.40 2.44 ;
        RECT  11.24 1.40 11.40 2.44 ;
        RECT  9.52 2.36 10.68 2.52 ;
    END
END MUX5SP4V1_0

MACRO MUX5SP2V1_0
    CLASS CORE ;
    FOREIGN MUX5SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 20.10  LAYER ME1  ;
        ANTENNADIFFAREA 8.51  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.42  LAYER ME1  ;
        ANTENNAMAXAREACAR 48.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.56 1.84 11.88 2.12 ;
        RECT  11.72 0.94 11.88 2.12 ;
        RECT  11.56 0.94 11.88 1.22 ;
        END
    END OUT
    PIN S2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.68 1.38 11.08 1.68 ;
        END
    END S2
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.60 1.26 7.88 1.68 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.46 0.50 1.74 ;
        END
    END S0
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.08 1.26 8.36 1.68 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.33  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 19.73  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.66 0.76 3.94 2.20 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.96  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 14.21  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.76 1.46 3.14 1.74 ;
        RECT  2.62 1.92 2.92 2.20 ;
        RECT  2.76 0.76 2.92 2.20 ;
        RECT  2.62 0.76 2.92 1.04 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.49  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 22.12  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.14 1.92 2.42 2.20 ;
        RECT  2.14 0.76 2.42 1.04 ;
        RECT  2.14 0.76 2.34 2.20 ;
        RECT  2.06 1.46 2.34 1.74 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.14  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.02  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.22 1.46 1.54 1.74 ;
        RECT  1.10 1.92 1.38 2.20 ;
        RECT  1.22 0.76 1.38 2.20 ;
        RECT  1.10 0.76 1.38 1.04 ;
        END
    END A
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 12.00 0.28 ;
        RECT  11.54 -0.28 11.82 0.32 ;
        RECT  11.04 0.94 11.32 1.22 ;
        RECT  11.10 -0.28 11.26 1.22 ;
        RECT  7.78 0.82 8.06 1.10 ;
        RECT  7.84 -0.28 8.00 1.10 ;
        RECT  4.76 0.96 5.04 1.24 ;
        RECT  4.82 -0.28 4.98 1.24 ;
        RECT  0.10 0.96 0.38 1.24 ;
        RECT  0.16 -0.28 0.32 1.24 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 12.00 3.48 ;
        RECT  11.54 2.88 11.82 3.48 ;
        RECT  10.95 2.62 11.23 3.48 ;
        RECT  7.82 2.62 8.10 3.48 ;
        RECT  4.59 2.62 4.87 3.48 ;
        RECT  0.10 1.90 0.38 2.18 ;
        RECT  0.16 1.90 0.32 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.96 0.90 1.24 ;
        RECT  0.68 1.40 1.04 1.68 ;
        RECT  0.68 0.96 0.84 2.18 ;
        RECT  0.62 1.90 0.90 2.18 ;
        RECT  3.30 0.44 4.38 0.60 ;
        RECT  4.10 0.44 4.38 0.72 ;
        RECT  3.14 0.76 3.46 1.04 ;
        RECT  3.30 0.44 3.46 2.20 ;
        RECT  3.14 1.92 3.46 2.20 ;
        RECT  1.62 0.76 1.90 1.04 ;
        RECT  1.70 0.76 1.86 2.20 ;
        RECT  1.62 1.92 1.90 2.20 ;
        RECT  1.74 1.92 1.90 2.52 ;
        RECT  1.74 2.36 4.44 2.52 ;
        RECT  4.16 2.28 4.44 2.56 ;
        RECT  5.32 0.76 5.60 1.04 ;
        RECT  5.38 0.76 5.54 2.20 ;
        RECT  5.32 1.92 5.60 2.20 ;
        RECT  6.34 0.76 6.64 1.04 ;
        RECT  4.24 0.96 4.52 1.24 ;
        RECT  4.30 0.96 4.46 2.12 ;
        RECT  6.34 0.76 6.50 2.20 ;
        RECT  4.24 1.84 4.52 2.12 ;
        RECT  4.24 1.96 5.16 2.12 ;
        RECT  6.34 1.92 6.64 2.20 ;
        RECT  5.00 1.96 5.16 2.52 ;
        RECT  6.36 1.92 6.52 2.52 ;
        RECT  5.00 2.36 6.52 2.52 ;
        RECT  7.26 0.82 7.54 1.10 ;
        RECT  7.12 1.40 7.42 1.68 ;
        RECT  7.26 0.82 7.42 2.12 ;
        RECT  7.26 1.84 7.54 2.12 ;
        RECT  5.96 0.44 6.96 0.60 ;
        RECT  5.96 0.44 6.12 1.04 ;
        RECT  5.84 0.76 6.12 1.04 ;
        RECT  8.88 0.76 9.16 1.04 ;
        RECT  5.90 0.76 6.06 2.20 ;
        RECT  8.94 0.76 9.10 2.20 ;
        RECT  5.84 1.92 6.12 2.20 ;
        RECT  8.88 1.92 9.16 2.20 ;
        RECT  6.80 0.44 6.96 2.44 ;
        RECT  8.88 1.92 9.04 2.44 ;
        RECT  6.80 2.28 9.04 2.44 ;
        RECT  8.52 0.44 10.08 0.60 ;
        RECT  9.92 0.76 10.20 1.04 ;
        RECT  8.30 0.82 8.68 1.10 ;
        RECT  9.92 0.44 10.08 2.20 ;
        RECT  8.52 0.44 8.68 2.12 ;
        RECT  8.30 1.84 8.68 2.12 ;
        RECT  9.92 1.92 10.20 2.20 ;
        RECT  10.36 0.94 10.80 1.22 ;
        RECT  10.24 1.40 10.52 1.68 ;
        RECT  10.36 0.94 10.52 2.12 ;
        RECT  10.36 1.84 10.80 2.12 ;
        RECT  9.40 0.76 9.68 1.04 ;
        RECT  11.24 1.40 11.56 1.68 ;
        RECT  9.46 0.76 9.62 2.20 ;
        RECT  9.40 1.92 9.68 2.20 ;
        RECT  9.52 1.92 9.68 2.52 ;
        RECT  10.52 2.28 11.40 2.44 ;
        RECT  11.24 1.40 11.40 2.44 ;
        RECT  9.52 2.36 10.68 2.52 ;
    END
END MUX5SP2V1_0

MACRO MUX5SP1V1_0
    CLASS CORE ;
    FOREIGN MUX5SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.14  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.02  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.22 1.46 1.54 1.74 ;
        RECT  1.10 1.92 1.38 2.20 ;
        RECT  1.22 0.76 1.38 2.20 ;
        RECT  1.10 0.76 1.38 1.04 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.49  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 22.12  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.14 1.92 2.42 2.20 ;
        RECT  2.14 0.76 2.42 1.04 ;
        RECT  2.14 0.76 2.34 2.20 ;
        RECT  2.06 1.46 2.34 1.74 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.96  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 14.21  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.76 1.46 3.14 1.74 ;
        RECT  2.62 1.92 2.92 2.20 ;
        RECT  2.76 0.76 2.92 2.20 ;
        RECT  2.62 0.76 2.92 1.04 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.33  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 19.73  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.66 0.76 3.94 2.20 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.08 1.26 8.36 1.68 ;
        END
    END E
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.46 0.50 1.74 ;
        END
    END S0
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.60 1.26 7.88 1.68 ;
        END
    END S1
    PIN S2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.77 1.40 11.19 1.68 ;
        END
    END S2
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 19.97  LAYER ME1  ;
        ANTENNADIFFAREA 8.13  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.34  LAYER ME1  ;
        ANTENNAMAXAREACAR 59.44  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.54 1.84 11.88 2.12 ;
        RECT  11.72 0.96 11.88 2.12 ;
        RECT  11.54 0.96 11.88 1.24 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 12.00 3.48 ;
        RECT  11.54 2.88 11.82 3.48 ;
        RECT  10.93 2.62 11.21 3.48 ;
        RECT  7.82 2.62 8.10 3.48 ;
        RECT  4.59 2.62 4.87 3.48 ;
        RECT  0.10 1.90 0.38 2.18 ;
        RECT  0.16 1.90 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 12.00 0.28 ;
        RECT  11.54 -0.28 11.82 0.32 ;
        RECT  11.02 0.96 11.30 1.24 ;
        RECT  11.08 -0.28 11.24 1.24 ;
        RECT  7.78 0.82 8.06 1.10 ;
        RECT  7.84 -0.28 8.00 1.10 ;
        RECT  4.76 0.96 5.04 1.24 ;
        RECT  4.82 -0.28 4.98 1.24 ;
        RECT  0.10 0.96 0.38 1.24 ;
        RECT  0.16 -0.28 0.32 1.24 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.96 0.90 1.24 ;
        RECT  0.68 1.40 1.04 1.68 ;
        RECT  0.68 0.96 0.84 2.18 ;
        RECT  0.62 1.90 0.90 2.18 ;
        RECT  3.30 0.44 4.38 0.60 ;
        RECT  4.10 0.44 4.38 0.72 ;
        RECT  3.14 0.76 3.46 1.04 ;
        RECT  3.30 0.44 3.46 2.20 ;
        RECT  3.14 1.92 3.46 2.20 ;
        RECT  1.62 0.76 1.90 1.04 ;
        RECT  1.70 0.76 1.86 2.20 ;
        RECT  1.62 1.92 1.90 2.20 ;
        RECT  1.74 1.92 1.90 2.52 ;
        RECT  1.74 2.36 4.44 2.52 ;
        RECT  4.16 2.28 4.44 2.56 ;
        RECT  5.32 0.76 5.60 1.04 ;
        RECT  5.38 0.76 5.54 2.20 ;
        RECT  5.32 1.92 5.60 2.20 ;
        RECT  6.34 0.76 6.64 1.04 ;
        RECT  4.24 0.96 4.52 1.24 ;
        RECT  4.30 0.96 4.46 2.12 ;
        RECT  6.34 0.76 6.50 2.20 ;
        RECT  4.24 1.84 4.52 2.12 ;
        RECT  4.24 1.96 5.16 2.12 ;
        RECT  6.34 1.92 6.64 2.20 ;
        RECT  5.00 1.96 5.16 2.52 ;
        RECT  6.36 1.92 6.52 2.52 ;
        RECT  5.00 2.36 6.52 2.52 ;
        RECT  7.26 0.82 7.54 1.10 ;
        RECT  7.12 1.40 7.42 1.68 ;
        RECT  7.26 0.82 7.42 2.12 ;
        RECT  7.26 1.84 7.54 2.12 ;
        RECT  5.96 0.44 6.96 0.60 ;
        RECT  5.96 0.44 6.12 1.04 ;
        RECT  5.84 0.76 6.12 1.04 ;
        RECT  8.88 0.76 9.16 1.04 ;
        RECT  5.90 0.76 6.06 2.20 ;
        RECT  8.94 0.76 9.10 2.20 ;
        RECT  5.84 1.92 6.12 2.20 ;
        RECT  8.88 1.92 9.16 2.20 ;
        RECT  6.80 0.44 6.96 2.44 ;
        RECT  8.88 1.92 9.04 2.44 ;
        RECT  6.80 2.28 9.04 2.44 ;
        RECT  8.52 0.44 10.08 0.60 ;
        RECT  9.92 0.76 10.20 1.04 ;
        RECT  8.30 0.82 8.68 1.10 ;
        RECT  9.92 0.44 10.08 2.20 ;
        RECT  8.52 0.44 8.68 2.12 ;
        RECT  8.30 1.84 8.68 2.12 ;
        RECT  9.92 1.92 10.20 2.20 ;
        RECT  10.36 0.96 10.78 1.24 ;
        RECT  10.24 1.40 10.52 1.68 ;
        RECT  10.36 0.96 10.52 2.12 ;
        RECT  10.36 1.84 10.78 2.12 ;
        RECT  9.40 0.76 9.68 1.04 ;
        RECT  9.46 0.76 9.62 2.20 ;
        RECT  9.40 1.92 9.68 2.20 ;
        RECT  9.52 1.92 9.68 2.52 ;
        RECT  10.52 2.28 11.64 2.44 ;
        RECT  9.52 2.36 10.68 2.52 ;
        RECT  11.36 2.28 11.64 2.56 ;
    END
END MUX5SP1V1_0

MACRO MUX4SP8V1_0
    CLASS CORE ;
    FOREIGN MUX4SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 16.83  LAYER ME1  ;
        ANTENNADIFFAREA 8.22  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.85  LAYER ME1  ;
        ANTENNAMAXAREACAR 19.69  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.40 1.84 9.68 2.12 ;
        RECT  9.40 0.96 9.68 1.24 ;
        RECT  9.40 0.96 9.56 2.12 ;
        RECT  8.52 1.52 9.56 1.68 ;
        RECT  8.36 1.84 8.68 2.12 ;
        RECT  8.52 0.96 8.68 2.12 ;
        RECT  8.36 0.96 8.68 1.24 ;
        END
    END OUT
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.56 1.38 7.88 1.70 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.40 0.50 1.68 ;
        END
    END S0
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.14  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 16.98  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.66 1.92 3.94 2.20 ;
        RECT  3.66 0.76 3.94 1.04 ;
        RECT  3.72 0.76 3.88 2.20 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.17  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.36  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.62 1.92 2.90 2.20 ;
        RECT  2.62 0.76 2.90 1.04 ;
        RECT  2.68 0.76 2.84 2.20 ;
        RECT  2.52 1.52 2.84 1.68 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.40  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 20.90  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.12 1.92 2.42 2.20 ;
        RECT  2.12 0.76 2.42 1.04 ;
        RECT  2.12 0.76 2.28 2.20 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.42  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 21.19  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.20 1.52 1.48 1.68 ;
        RECT  1.10 1.92 1.38 2.20 ;
        RECT  1.10 0.76 1.38 1.04 ;
        RECT  1.20 0.76 1.36 2.20 ;
        END
    END A
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 10.40 0.28 ;
        RECT  9.94 -0.28 10.22 0.32 ;
        RECT  9.92 0.56 10.20 0.84 ;
        RECT  9.98 -0.28 10.14 0.84 ;
        RECT  8.88 0.56 9.16 0.84 ;
        RECT  8.94 -0.28 9.10 0.84 ;
        RECT  7.84 0.94 8.12 1.22 ;
        RECT  7.90 -0.28 8.06 1.22 ;
        RECT  4.76 0.96 5.04 1.24 ;
        RECT  4.82 -0.28 4.98 1.24 ;
        RECT  0.10 0.96 0.38 1.24 ;
        RECT  0.16 -0.28 0.32 1.24 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 10.40 3.48 ;
        RECT  9.94 2.88 10.22 3.48 ;
        RECT  9.92 2.24 10.20 2.52 ;
        RECT  9.98 2.24 10.14 3.48 ;
        RECT  8.88 2.24 9.16 2.52 ;
        RECT  8.94 2.24 9.10 3.48 ;
        RECT  7.75 2.62 8.03 3.48 ;
        RECT  4.59 2.62 4.87 3.48 ;
        RECT  0.10 1.84 0.38 2.12 ;
        RECT  0.16 1.84 0.32 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.96 0.90 1.24 ;
        RECT  0.72 1.40 1.04 1.68 ;
        RECT  0.72 0.96 0.88 2.12 ;
        RECT  0.62 1.84 0.90 2.12 ;
        RECT  3.20 0.44 4.38 0.60 ;
        RECT  4.10 0.44 4.38 0.72 ;
        RECT  3.14 0.76 3.42 1.04 ;
        RECT  3.20 0.44 3.36 2.20 ;
        RECT  3.14 1.92 3.42 2.20 ;
        RECT  1.62 0.76 1.90 1.04 ;
        RECT  1.62 1.92 1.90 2.20 ;
        RECT  1.68 0.76 1.84 2.52 ;
        RECT  1.68 2.36 4.44 2.52 ;
        RECT  4.16 2.28 4.44 2.56 ;
        RECT  5.32 0.76 5.60 1.04 ;
        RECT  5.38 0.76 5.54 2.20 ;
        RECT  5.32 1.92 5.60 2.20 ;
        RECT  6.36 0.76 6.64 1.04 ;
        RECT  4.24 0.96 4.52 1.24 ;
        RECT  4.30 0.96 4.46 2.12 ;
        RECT  6.38 0.76 6.54 2.20 ;
        RECT  4.24 1.84 4.52 2.12 ;
        RECT  4.24 1.96 5.16 2.12 ;
        RECT  6.36 1.92 6.64 2.20 ;
        RECT  5.00 1.96 5.16 2.52 ;
        RECT  6.36 1.92 6.52 2.52 ;
        RECT  5.00 2.36 6.52 2.52 ;
        RECT  7.24 0.94 7.60 1.22 ;
        RECT  7.12 1.40 7.40 1.68 ;
        RECT  7.24 0.94 7.40 2.14 ;
        RECT  7.24 1.86 7.60 2.14 ;
        RECT  5.96 0.44 6.96 0.60 ;
        RECT  5.96 0.44 6.12 1.04 ;
        RECT  5.84 0.76 6.12 1.04 ;
        RECT  8.04 1.40 8.36 1.68 ;
        RECT  5.90 0.76 6.06 2.20 ;
        RECT  5.84 1.92 6.12 2.20 ;
        RECT  6.80 0.44 6.96 2.46 ;
        RECT  8.04 1.40 8.20 2.46 ;
        RECT  6.80 2.30 8.20 2.46 ;
    END
END MUX4SP8V1_0

MACRO MUX4SP4V1_0
    CLASS CORE ;
    FOREIGN MUX4SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.42  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 21.19  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.20 1.52 1.48 1.68 ;
        RECT  1.10 1.92 1.38 2.20 ;
        RECT  1.10 0.76 1.38 1.04 ;
        RECT  1.20 0.76 1.36 2.20 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.12  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 16.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.12 1.92 2.42 2.20 ;
        RECT  2.12 0.76 2.42 1.04 ;
        RECT  2.12 0.76 2.28 2.20 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.17  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.36  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.62 1.92 2.90 2.20 ;
        RECT  2.62 0.76 2.90 1.04 ;
        RECT  2.68 0.76 2.84 2.20 ;
        RECT  2.52 1.52 2.84 1.68 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.87  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 12.93  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.66 1.92 3.94 2.20 ;
        RECT  3.66 0.76 3.94 1.04 ;
        RECT  3.72 0.76 3.88 2.20 ;
        END
    END D
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.40 0.50 1.68 ;
        END
    END S0
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.56 1.36 7.88 1.68 ;
        END
    END S1
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 15.05  LAYER ME1  ;
        ANTENNADIFFAREA 6.52  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER ME1  ;
        ANTENNAMAXAREACAR 30.73  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.36 1.84 8.68 2.12 ;
        RECT  8.52 0.92 8.68 2.12 ;
        RECT  8.36 0.92 8.68 1.20 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 9.60 3.48 ;
        RECT  8.94 2.88 9.42 3.48 ;
        RECT  8.88 2.16 9.16 2.44 ;
        RECT  8.94 2.16 9.10 3.48 ;
        RECT  7.75 2.62 8.03 3.48 ;
        RECT  4.59 2.62 4.87 3.48 ;
        RECT  0.10 1.84 0.38 2.12 ;
        RECT  0.16 1.84 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 9.60 0.28 ;
        RECT  8.94 -0.28 9.42 0.32 ;
        RECT  8.88 0.60 9.16 0.88 ;
        RECT  8.94 -0.28 9.10 0.88 ;
        RECT  7.84 0.92 8.12 1.20 ;
        RECT  7.90 -0.28 8.06 1.20 ;
        RECT  4.76 0.96 5.04 1.24 ;
        RECT  4.82 -0.28 4.98 1.24 ;
        RECT  0.10 0.96 0.38 1.24 ;
        RECT  0.16 -0.28 0.32 1.24 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.96 0.90 1.24 ;
        RECT  0.72 1.40 1.04 1.68 ;
        RECT  0.72 0.96 0.88 2.12 ;
        RECT  0.62 1.84 0.90 2.12 ;
        RECT  3.20 0.44 4.38 0.60 ;
        RECT  4.10 0.44 4.38 0.72 ;
        RECT  3.14 0.76 3.42 1.04 ;
        RECT  3.20 0.44 3.36 2.20 ;
        RECT  3.14 1.92 3.42 2.20 ;
        RECT  1.62 0.76 1.90 1.04 ;
        RECT  1.62 1.92 1.90 2.20 ;
        RECT  1.68 0.76 1.84 2.52 ;
        RECT  1.68 2.36 4.44 2.52 ;
        RECT  4.16 2.28 4.44 2.56 ;
        RECT  5.32 0.76 5.60 1.04 ;
        RECT  5.38 0.76 5.54 2.20 ;
        RECT  5.32 1.92 5.60 2.20 ;
        RECT  6.36 0.76 6.64 1.04 ;
        RECT  4.24 0.96 4.52 1.24 ;
        RECT  4.30 0.96 4.46 2.12 ;
        RECT  6.38 0.76 6.54 2.20 ;
        RECT  4.24 1.84 4.52 2.12 ;
        RECT  4.24 1.96 5.16 2.12 ;
        RECT  6.36 1.92 6.64 2.20 ;
        RECT  5.00 1.96 5.16 2.52 ;
        RECT  6.36 1.92 6.52 2.52 ;
        RECT  5.00 2.36 6.52 2.52 ;
        RECT  7.24 0.92 7.60 1.20 ;
        RECT  7.12 1.40 7.40 1.68 ;
        RECT  7.24 0.92 7.40 2.12 ;
        RECT  7.24 1.84 7.60 2.12 ;
        RECT  5.96 0.44 6.96 0.60 ;
        RECT  5.96 0.44 6.12 1.04 ;
        RECT  5.84 0.76 6.12 1.04 ;
        RECT  8.04 1.40 8.36 1.68 ;
        RECT  5.90 0.76 6.06 2.20 ;
        RECT  5.84 1.92 6.12 2.20 ;
        RECT  6.80 0.44 6.96 2.44 ;
        RECT  8.04 1.40 8.20 2.44 ;
        RECT  6.80 2.28 8.20 2.44 ;
    END
END MUX4SP4V1_0

MACRO MUX4SP2V1_0
    CLASS CORE ;
    FOREIGN MUX4SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 13.86  LAYER ME1  ;
        ANTENNADIFFAREA 5.79  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.35  LAYER ME1  ;
        ANTENNAMAXAREACAR 40.11  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.36 1.84 8.68 2.12 ;
        RECT  8.52 0.92 8.68 2.12 ;
        RECT  8.36 0.92 8.68 1.20 ;
        END
    END OUT
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.56 1.36 7.88 1.68 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.40 0.50 1.68 ;
        END
    END S0
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.14  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 16.98  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.66 1.92 3.94 2.20 ;
        RECT  3.66 0.76 3.94 1.04 ;
        RECT  3.72 0.76 3.88 2.20 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.17  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.36  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.62 1.92 2.90 2.20 ;
        RECT  2.62 0.76 2.90 1.04 ;
        RECT  2.68 0.76 2.84 2.20 ;
        RECT  2.52 1.52 2.84 1.68 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.40  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 20.90  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.12 1.92 2.42 2.20 ;
        RECT  2.12 0.76 2.42 1.04 ;
        RECT  2.12 0.76 2.28 2.20 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.42  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 21.19  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.20 1.52 1.48 1.68 ;
        RECT  1.10 1.92 1.38 2.20 ;
        RECT  1.10 0.76 1.38 1.04 ;
        RECT  1.20 0.76 1.36 2.20 ;
        END
    END A
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 8.80 0.28 ;
        RECT  8.34 -0.28 8.62 0.32 ;
        RECT  7.84 0.92 8.12 1.20 ;
        RECT  7.90 -0.28 8.06 1.20 ;
        RECT  4.76 0.96 5.04 1.24 ;
        RECT  4.82 -0.28 4.98 1.24 ;
        RECT  0.10 0.96 0.38 1.24 ;
        RECT  0.16 -0.28 0.32 1.24 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 8.80 3.48 ;
        RECT  8.34 2.88 8.62 3.48 ;
        RECT  7.75 2.62 8.03 3.48 ;
        RECT  4.59 2.62 4.87 3.48 ;
        RECT  0.10 1.84 0.38 2.12 ;
        RECT  0.16 1.84 0.32 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.96 0.90 1.24 ;
        RECT  0.72 1.40 1.04 1.68 ;
        RECT  0.72 0.96 0.88 2.12 ;
        RECT  0.62 1.84 0.90 2.12 ;
        RECT  3.20 0.44 4.38 0.60 ;
        RECT  4.10 0.44 4.38 0.72 ;
        RECT  3.14 0.76 3.42 1.04 ;
        RECT  3.20 0.44 3.36 2.20 ;
        RECT  3.14 1.92 3.42 2.20 ;
        RECT  1.62 0.76 1.90 1.04 ;
        RECT  1.62 1.92 1.90 2.20 ;
        RECT  1.68 0.76 1.84 2.52 ;
        RECT  1.68 2.36 4.44 2.52 ;
        RECT  4.16 2.28 4.44 2.56 ;
        RECT  5.32 0.76 5.60 1.04 ;
        RECT  5.38 0.76 5.54 2.20 ;
        RECT  5.32 1.92 5.60 2.20 ;
        RECT  6.36 0.76 6.64 1.04 ;
        RECT  4.24 0.96 4.52 1.24 ;
        RECT  4.30 0.96 4.46 2.12 ;
        RECT  6.38 0.76 6.54 2.20 ;
        RECT  4.24 1.84 4.52 2.12 ;
        RECT  4.24 1.96 5.16 2.12 ;
        RECT  6.36 1.92 6.64 2.20 ;
        RECT  5.00 1.96 5.16 2.52 ;
        RECT  6.36 1.92 6.52 2.52 ;
        RECT  5.00 2.36 6.52 2.52 ;
        RECT  7.24 0.92 7.60 1.20 ;
        RECT  7.12 1.40 7.40 1.68 ;
        RECT  7.24 0.92 7.40 2.12 ;
        RECT  7.24 1.84 7.60 2.12 ;
        RECT  5.96 0.44 6.96 0.60 ;
        RECT  5.96 0.44 6.12 1.04 ;
        RECT  5.84 0.76 6.12 1.04 ;
        RECT  8.04 1.40 8.36 1.68 ;
        RECT  5.90 0.76 6.06 2.20 ;
        RECT  5.84 1.92 6.12 2.20 ;
        RECT  6.80 0.44 6.96 2.44 ;
        RECT  8.04 1.40 8.20 2.44 ;
        RECT  6.80 2.28 8.20 2.44 ;
    END
END MUX4SP2V1_0

MACRO MUX4SP1V1_0
    CLASS CORE ;
    FOREIGN MUX4SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.42  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 21.19  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.20 1.52 1.48 1.68 ;
        RECT  1.10 1.92 1.38 2.20 ;
        RECT  1.10 0.76 1.38 1.04 ;
        RECT  1.20 0.76 1.36 2.20 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.12  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 16.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.12 1.92 2.42 2.20 ;
        RECT  2.12 0.76 2.42 1.04 ;
        RECT  2.12 0.76 2.28 2.20 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.17  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.36  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.62 1.92 2.90 2.20 ;
        RECT  2.62 0.76 2.90 1.04 ;
        RECT  2.68 0.76 2.84 2.20 ;
        RECT  2.52 1.52 2.84 1.68 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.87  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 12.93  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.66 1.92 3.94 2.20 ;
        RECT  3.66 0.76 3.94 1.04 ;
        RECT  3.72 0.76 3.88 2.20 ;
        END
    END D
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.40 0.50 1.68 ;
        END
    END S0
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.58 1.40 8.00 1.68 ;
        END
    END S1
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 14.01  LAYER ME1  ;
        ANTENNADIFFAREA 5.43  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.27  LAYER ME1  ;
        ANTENNAMAXAREACAR 52.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.30 1.84 8.68 2.12 ;
        RECT  8.52 0.96 8.68 2.12 ;
        RECT  8.30 0.96 8.68 1.24 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 8.80 3.48 ;
        RECT  8.34 2.88 8.62 3.48 ;
        RECT  7.69 2.62 7.97 3.48 ;
        RECT  4.59 2.62 4.87 3.48 ;
        RECT  0.10 1.84 0.38 2.12 ;
        RECT  0.16 1.84 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 8.80 0.28 ;
        RECT  8.34 -0.28 8.62 0.32 ;
        RECT  7.78 0.96 8.06 1.24 ;
        RECT  7.84 -0.28 8.00 1.24 ;
        RECT  4.76 0.96 5.04 1.24 ;
        RECT  4.82 -0.28 4.98 1.24 ;
        RECT  0.10 0.96 0.38 1.24 ;
        RECT  0.16 -0.28 0.32 1.24 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.96 0.90 1.24 ;
        RECT  0.72 1.40 1.04 1.68 ;
        RECT  0.72 0.96 0.88 2.12 ;
        RECT  0.62 1.84 0.90 2.12 ;
        RECT  3.20 0.44 4.38 0.60 ;
        RECT  4.10 0.44 4.38 0.72 ;
        RECT  3.14 0.76 3.42 1.04 ;
        RECT  3.20 0.44 3.36 2.20 ;
        RECT  3.14 1.92 3.42 2.20 ;
        RECT  1.62 0.76 1.90 1.04 ;
        RECT  1.62 1.92 1.90 2.20 ;
        RECT  1.68 0.76 1.84 2.52 ;
        RECT  1.68 2.36 4.44 2.52 ;
        RECT  4.16 2.28 4.44 2.56 ;
        RECT  5.32 0.76 5.60 1.04 ;
        RECT  5.38 0.76 5.54 2.20 ;
        RECT  5.32 1.92 5.60 2.20 ;
        RECT  6.36 0.76 6.64 1.04 ;
        RECT  4.24 0.96 4.52 1.24 ;
        RECT  4.30 0.96 4.46 2.12 ;
        RECT  6.38 0.76 6.54 2.20 ;
        RECT  4.24 1.84 4.52 2.12 ;
        RECT  4.24 1.96 5.16 2.12 ;
        RECT  6.36 1.92 6.64 2.20 ;
        RECT  5.00 1.96 5.16 2.52 ;
        RECT  6.36 1.92 6.52 2.52 ;
        RECT  5.00 2.36 6.52 2.52 ;
        RECT  7.26 0.96 7.54 1.24 ;
        RECT  7.12 1.40 7.42 1.68 ;
        RECT  7.26 0.96 7.42 2.12 ;
        RECT  7.26 1.84 7.54 2.12 ;
        RECT  5.96 0.44 6.96 0.60 ;
        RECT  5.96 0.44 6.12 1.04 ;
        RECT  5.84 0.76 6.12 1.04 ;
        RECT  5.90 0.76 6.06 2.20 ;
        RECT  5.84 1.92 6.12 2.20 ;
        RECT  6.80 0.44 6.96 2.44 ;
        RECT  6.80 2.28 8.40 2.44 ;
        RECT  8.12 2.28 8.40 2.56 ;
    END
END MUX4SP1V1_0

MACRO MUX4LSP8V1_0
    CLASS CORE ;
    FOREIGN MUX4LSP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 13.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 21.74  LAYER ME1  ;
        ANTENNADIFFAREA 11.52  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.87  LAYER ME1  ;
        ANTENNAMAXAREACAR 24.89  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.00 1.84 12.28 2.12 ;
        RECT  8.88 1.08 12.28 1.24 ;
        RECT  12.00 0.96 12.28 1.24 ;
        RECT  10.96 1.84 12.28 2.00 ;
        RECT  11.72 1.08 11.88 2.00 ;
        RECT  10.96 1.84 11.24 2.12 ;
        RECT  10.96 0.96 11.24 1.24 ;
        RECT  9.92 0.96 10.20 1.24 ;
        RECT  8.88 0.96 9.16 1.24 ;
        END
    END OUT
    PIN EN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.73 1.40 11.15 1.68 ;
        END
    END EN
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.60 1.26 7.88 1.68 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.40 0.50 1.68 ;
        END
    END S0
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.84  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 12.57  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.66 1.92 3.94 2.20 ;
        RECT  3.66 0.76 3.94 1.04 ;
        RECT  3.72 0.76 3.88 2.20 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.17  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.38  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.76 1.52 3.08 1.68 ;
        RECT  2.62 1.92 2.92 2.20 ;
        RECT  2.76 0.76 2.92 2.20 ;
        RECT  2.62 0.76 2.92 1.04 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.39  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 20.74  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.12 1.92 2.42 2.20 ;
        RECT  2.12 0.76 2.42 1.04 ;
        RECT  2.12 0.76 2.28 2.20 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.41  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 20.98  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.22 1.52 1.48 1.68 ;
        RECT  1.10 1.92 1.38 2.20 ;
        RECT  1.22 0.76 1.38 2.20 ;
        RECT  1.10 0.76 1.38 1.04 ;
        END
    END A
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 13.20 0.28 ;
        RECT  12.58 -0.28 13.02 0.32 ;
        RECT  12.52 0.54 12.80 0.82 ;
        RECT  12.58 -0.28 12.74 0.82 ;
        RECT  11.48 0.54 11.76 0.82 ;
        RECT  11.54 -0.28 11.70 0.82 ;
        RECT  10.44 0.54 10.72 0.82 ;
        RECT  10.50 -0.28 10.66 0.82 ;
        RECT  9.40 0.54 9.68 0.82 ;
        RECT  9.46 -0.28 9.62 0.82 ;
        RECT  8.36 0.54 8.64 0.82 ;
        RECT  8.42 -0.28 8.58 0.82 ;
        RECT  7.78 0.82 8.06 1.10 ;
        RECT  7.84 -0.28 8.00 1.10 ;
        RECT  4.76 0.96 5.04 1.24 ;
        RECT  4.82 -0.28 4.98 1.24 ;
        RECT  0.10 0.96 0.38 1.24 ;
        RECT  0.16 -0.28 0.32 1.24 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 13.20 3.48 ;
        RECT  12.74 2.88 13.02 3.48 ;
        RECT  9.92 2.26 10.20 2.54 ;
        RECT  9.98 2.26 10.14 3.48 ;
        RECT  8.88 2.26 9.16 2.54 ;
        RECT  8.94 2.26 9.10 3.48 ;
        RECT  7.82 2.62 8.10 3.48 ;
        RECT  4.58 2.62 4.86 3.48 ;
        RECT  0.10 1.84 0.38 2.12 ;
        RECT  0.16 1.84 0.32 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.96 0.90 1.24 ;
        RECT  0.68 1.40 1.04 1.68 ;
        RECT  0.68 0.96 0.84 2.12 ;
        RECT  0.62 1.84 0.90 2.12 ;
        RECT  3.26 0.44 4.38 0.60 ;
        RECT  4.10 0.44 4.38 0.72 ;
        RECT  3.26 0.44 3.42 1.04 ;
        RECT  3.14 0.76 3.42 1.04 ;
        RECT  3.24 0.76 3.40 2.20 ;
        RECT  3.14 1.92 3.42 2.20 ;
        RECT  1.62 0.76 1.90 1.04 ;
        RECT  1.68 0.76 1.84 2.20 ;
        RECT  1.62 1.92 1.90 2.20 ;
        RECT  1.74 1.92 1.90 2.52 ;
        RECT  1.74 2.36 4.43 2.52 ;
        RECT  4.15 2.28 4.43 2.56 ;
        RECT  5.32 0.76 5.60 1.04 ;
        RECT  5.38 0.76 5.54 2.20 ;
        RECT  5.32 1.92 5.60 2.20 ;
        RECT  6.36 0.76 6.64 1.04 ;
        RECT  4.24 0.96 4.52 1.24 ;
        RECT  4.30 0.96 4.46 2.12 ;
        RECT  6.38 0.76 6.54 2.20 ;
        RECT  4.24 1.84 4.52 2.12 ;
        RECT  4.24 1.96 5.16 2.12 ;
        RECT  6.36 1.92 6.64 2.20 ;
        RECT  5.00 1.96 5.16 2.53 ;
        RECT  6.36 1.92 6.52 2.53 ;
        RECT  5.00 2.37 6.52 2.53 ;
        RECT  7.26 0.82 7.54 1.10 ;
        RECT  7.12 1.40 7.42 1.68 ;
        RECT  7.26 0.82 7.42 2.12 ;
        RECT  7.26 1.84 7.54 2.12 ;
        RECT  5.96 0.44 6.96 0.60 ;
        RECT  5.96 0.44 6.12 1.04 ;
        RECT  5.84 0.76 6.12 1.04 ;
        RECT  8.04 1.46 8.94 1.62 ;
        RECT  8.66 1.40 8.94 1.68 ;
        RECT  5.90 0.76 6.06 2.20 ;
        RECT  5.84 1.92 6.12 2.20 ;
        RECT  6.80 0.44 6.96 2.44 ;
        RECT  8.04 1.46 8.20 2.44 ;
        RECT  6.80 2.28 8.20 2.44 ;
        RECT  8.36 1.84 10.72 2.00 ;
        RECT  8.36 1.84 8.64 2.12 ;
        RECT  9.40 1.84 9.68 2.12 ;
        RECT  10.44 1.84 10.72 2.12 ;
        RECT  10.56 1.84 10.72 2.54 ;
        RECT  11.48 2.26 11.76 2.54 ;
        RECT  12.52 2.26 12.80 2.54 ;
        RECT  10.56 2.38 12.80 2.54 ;
    END
END MUX4LSP8V1_0

MACRO MUX4LSP4V1_0
    CLASS CORE ;
    FOREIGN MUX4LSP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 18.20  LAYER ME1  ;
        ANTENNADIFFAREA 8.41  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.51  LAYER ME1  ;
        ANTENNAMAXAREACAR 35.77  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.92 1.84 10.28 2.12 ;
        RECT  10.12 0.96 10.28 2.12 ;
        RECT  8.88 1.08 10.28 1.24 ;
        RECT  9.92 0.96 10.28 1.24 ;
        RECT  8.88 0.96 9.16 1.24 ;
        END
    END OUT
    PIN EN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.31  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.52 1.40 9.94 1.68 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.41  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 20.98  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.22 1.52 1.48 1.68 ;
        RECT  1.10 1.92 1.38 2.20 ;
        RECT  1.22 0.76 1.38 2.20 ;
        RECT  1.10 0.76 1.38 1.04 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.10  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 16.38  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.12 1.92 2.42 2.20 ;
        RECT  2.12 0.76 2.42 1.04 ;
        RECT  2.12 0.76 2.28 2.20 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.17  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.38  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.76 1.52 3.08 1.68 ;
        RECT  2.62 1.92 2.92 2.20 ;
        RECT  2.76 0.76 2.92 2.20 ;
        RECT  2.62 0.76 2.92 1.04 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.87  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 12.95  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.66 1.92 3.94 2.20 ;
        RECT  3.66 0.76 3.94 1.04 ;
        RECT  3.72 0.76 3.88 2.20 ;
        END
    END D
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.40 0.50 1.68 ;
        END
    END S0
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.60 1.26 7.88 1.68 ;
        END
    END S1
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 11.20 0.28 ;
        RECT  10.50 -0.28 11.02 0.32 ;
        RECT  10.44 0.60 10.72 0.88 ;
        RECT  10.50 -0.28 10.66 0.88 ;
        RECT  9.40 0.60 9.68 0.88 ;
        RECT  9.46 -0.28 9.62 0.88 ;
        RECT  8.36 0.60 8.64 0.88 ;
        RECT  8.42 -0.28 8.58 0.88 ;
        RECT  7.78 0.82 8.06 1.10 ;
        RECT  7.84 -0.28 8.00 1.10 ;
        RECT  4.76 0.96 5.04 1.24 ;
        RECT  4.82 -0.28 4.98 1.24 ;
        RECT  0.10 0.96 0.38 1.24 ;
        RECT  0.16 -0.28 0.32 1.24 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 11.20 3.48 ;
        RECT  10.74 2.88 11.02 3.48 ;
        RECT  8.88 2.20 9.16 2.48 ;
        RECT  8.94 2.20 9.10 3.48 ;
        RECT  7.82 2.62 8.10 3.48 ;
        RECT  4.58 2.62 4.86 3.48 ;
        RECT  0.10 1.84 0.38 2.12 ;
        RECT  0.16 1.84 0.32 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.96 0.90 1.24 ;
        RECT  0.68 1.40 1.04 1.68 ;
        RECT  0.68 0.96 0.84 2.12 ;
        RECT  0.62 1.84 0.90 2.12 ;
        RECT  3.26 0.44 4.38 0.60 ;
        RECT  4.10 0.44 4.38 0.72 ;
        RECT  3.26 0.44 3.42 1.04 ;
        RECT  3.14 0.76 3.42 1.04 ;
        RECT  3.24 0.76 3.40 2.20 ;
        RECT  3.14 1.92 3.42 2.20 ;
        RECT  1.62 0.76 1.90 1.04 ;
        RECT  1.68 0.76 1.84 2.20 ;
        RECT  1.62 1.92 1.90 2.20 ;
        RECT  1.74 1.92 1.90 2.52 ;
        RECT  1.74 2.36 4.43 2.52 ;
        RECT  4.15 2.28 4.43 2.56 ;
        RECT  5.32 0.76 5.60 1.04 ;
        RECT  5.38 0.76 5.54 2.20 ;
        RECT  5.32 1.92 5.60 2.20 ;
        RECT  6.36 0.76 6.64 1.04 ;
        RECT  4.24 0.96 4.52 1.24 ;
        RECT  4.30 0.96 4.46 2.12 ;
        RECT  6.38 0.76 6.54 2.20 ;
        RECT  4.24 1.84 4.52 2.12 ;
        RECT  4.24 1.96 5.16 2.12 ;
        RECT  6.36 1.92 6.64 2.20 ;
        RECT  5.00 1.96 5.16 2.53 ;
        RECT  6.36 1.92 6.52 2.53 ;
        RECT  5.00 2.37 6.52 2.53 ;
        RECT  7.26 0.82 7.54 1.10 ;
        RECT  7.12 1.40 7.42 1.68 ;
        RECT  7.26 0.82 7.42 2.12 ;
        RECT  7.26 1.84 7.54 2.12 ;
        RECT  5.96 0.44 6.96 0.60 ;
        RECT  5.96 0.44 6.12 1.04 ;
        RECT  5.84 0.76 6.12 1.04 ;
        RECT  8.04 1.46 8.94 1.62 ;
        RECT  8.66 1.40 8.94 1.68 ;
        RECT  5.90 0.76 6.06 2.20 ;
        RECT  5.84 1.92 6.12 2.20 ;
        RECT  6.80 0.44 6.96 2.44 ;
        RECT  8.04 1.46 8.20 2.44 ;
        RECT  6.80 2.28 8.20 2.44 ;
        RECT  8.36 1.84 9.68 2.00 ;
        RECT  8.36 1.84 8.64 2.12 ;
        RECT  9.40 1.84 9.68 2.12 ;
        RECT  9.52 1.84 9.68 2.48 ;
        RECT  10.44 2.20 10.72 2.48 ;
        RECT  9.52 2.32 10.72 2.48 ;
    END
END MUX4LSP4V1_0

MACRO MUX4LSP2V1_0
    CLASS CORE ;
    FOREIGN MUX4LSP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 15.29  LAYER ME1  ;
        ANTENNADIFFAREA 6.87  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.35  LAYER ME1  ;
        ANTENNAMAXAREACAR 43.64  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.86 1.96 9.48 2.12 ;
        RECT  9.32 1.08 9.48 2.12 ;
        RECT  8.34 1.08 9.48 1.24 ;
        RECT  8.86 1.84 9.14 2.12 ;
        RECT  8.34 0.96 8.62 1.24 ;
        END
    END OUT
    PIN EN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.15  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.72 1.40 9.14 1.68 ;
        END
    END EN
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.56 1.40 7.98 1.68 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.40 0.50 1.68 ;
        END
    END S0
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.84  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 12.57  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.66 1.92 3.94 2.20 ;
        RECT  3.66 0.76 3.94 1.04 ;
        RECT  3.72 0.76 3.88 2.20 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.17  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.38  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.76 1.52 3.08 1.68 ;
        RECT  2.62 1.92 2.92 2.20 ;
        RECT  2.76 0.76 2.92 2.20 ;
        RECT  2.62 0.76 2.92 1.04 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.39  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 20.74  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.12 1.92 2.42 2.20 ;
        RECT  2.12 0.76 2.42 1.04 ;
        RECT  2.12 0.76 2.28 2.20 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.41  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 20.98  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.22 1.52 1.48 1.68 ;
        RECT  1.10 1.92 1.38 2.20 ;
        RECT  1.22 0.76 1.38 2.20 ;
        RECT  1.10 0.76 1.38 1.04 ;
        END
    END A
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 9.60 3.48 ;
        RECT  9.14 2.88 9.42 3.48 ;
        RECT  7.78 2.62 8.06 3.48 ;
        RECT  4.58 2.62 4.86 3.48 ;
        RECT  0.10 1.84 0.38 2.12 ;
        RECT  0.16 1.84 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 9.60 0.28 ;
        RECT  8.92 -0.28 9.42 0.32 ;
        RECT  8.86 0.62 9.14 0.90 ;
        RECT  8.92 -0.28 9.08 0.90 ;
        RECT  7.82 0.62 8.10 0.90 ;
        RECT  7.88 -0.28 8.04 0.90 ;
        RECT  4.76 0.96 5.04 1.24 ;
        RECT  4.82 -0.28 4.98 1.24 ;
        RECT  0.10 0.96 0.38 1.24 ;
        RECT  0.16 -0.28 0.32 1.24 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.96 0.90 1.24 ;
        RECT  0.68 1.40 1.04 1.68 ;
        RECT  0.68 0.96 0.84 2.12 ;
        RECT  0.62 1.84 0.90 2.12 ;
        RECT  3.26 0.44 4.38 0.60 ;
        RECT  4.10 0.44 4.38 0.72 ;
        RECT  3.26 0.44 3.42 1.04 ;
        RECT  3.14 0.76 3.42 1.04 ;
        RECT  3.24 0.76 3.40 2.20 ;
        RECT  3.14 1.92 3.42 2.20 ;
        RECT  1.62 0.76 1.90 1.04 ;
        RECT  1.68 0.76 1.84 2.20 ;
        RECT  1.62 1.92 1.90 2.20 ;
        RECT  1.74 1.92 1.90 2.52 ;
        RECT  1.74 2.36 4.43 2.52 ;
        RECT  4.15 2.28 4.43 2.56 ;
        RECT  5.32 0.76 5.60 1.04 ;
        RECT  5.38 0.76 5.54 2.20 ;
        RECT  5.32 1.92 5.60 2.20 ;
        RECT  6.36 0.76 6.64 1.04 ;
        RECT  4.24 0.96 4.52 1.24 ;
        RECT  4.30 0.96 4.46 2.12 ;
        RECT  6.38 0.76 6.54 2.20 ;
        RECT  4.24 1.84 4.52 2.12 ;
        RECT  4.24 1.96 5.16 2.12 ;
        RECT  6.36 1.92 6.64 2.20 ;
        RECT  5.00 1.96 5.16 2.53 ;
        RECT  6.36 1.92 6.52 2.53 ;
        RECT  5.00 2.37 6.52 2.53 ;
        RECT  7.24 0.96 7.54 1.24 ;
        RECT  7.12 1.40 7.40 1.68 ;
        RECT  7.24 0.96 7.40 2.12 ;
        RECT  7.24 1.84 7.54 2.12 ;
        RECT  5.96 0.44 6.96 0.60 ;
        RECT  5.96 0.44 6.12 1.04 ;
        RECT  5.84 0.76 6.12 1.04 ;
        RECT  8.14 1.40 8.42 1.68 ;
        RECT  5.90 0.76 6.06 2.20 ;
        RECT  5.84 1.92 6.12 2.20 ;
        RECT  6.80 0.44 6.96 2.44 ;
        RECT  8.16 1.40 8.32 2.44 ;
        RECT  6.80 2.28 8.32 2.44 ;
    END
END MUX4LSP2V1_0

MACRO MUX4LSP1V1_0
    CLASS CORE ;
    FOREIGN MUX4LSP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.41  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 20.98  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.22 1.52 1.48 1.68 ;
        RECT  1.10 1.92 1.38 2.20 ;
        RECT  1.22 0.76 1.38 2.20 ;
        RECT  1.10 0.76 1.38 1.04 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.10  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 16.38  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.12 1.92 2.42 2.20 ;
        RECT  2.12 0.76 2.42 1.04 ;
        RECT  2.12 0.76 2.28 2.20 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.17  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.38  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.76 1.52 3.08 1.68 ;
        RECT  2.62 1.92 2.92 2.20 ;
        RECT  2.76 0.76 2.92 2.20 ;
        RECT  2.62 0.76 2.92 1.04 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.87  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 12.95  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.66 1.92 3.94 2.20 ;
        RECT  3.66 0.76 3.94 1.04 ;
        RECT  3.72 0.76 3.88 2.20 ;
        END
    END D
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.40 0.50 1.68 ;
        END
    END S0
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.60 1.26 7.88 1.68 ;
        END
    END S1
    PIN EN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.08 1.26 8.36 1.68 ;
        END
    END EN
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 15.22  LAYER ME1  ;
        ANTENNADIFFAREA 6.07  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.27  LAYER ME1  ;
        ANTENNAMAXAREACAR 56.63  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.82 1.84 9.10 2.12 ;
        RECT  8.92 1.02 9.08 2.12 ;
        RECT  8.50 1.02 9.08 1.18 ;
        RECT  8.50 0.54 8.66 1.18 ;
        RECT  8.30 0.54 8.66 0.82 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 9.60 3.48 ;
        RECT  9.14 2.88 9.42 3.48 ;
        RECT  7.82 2.62 8.10 3.48 ;
        RECT  4.58 2.62 4.86 3.48 ;
        RECT  0.10 1.84 0.38 2.12 ;
        RECT  0.16 1.84 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 9.60 0.28 ;
        RECT  8.88 -0.28 9.42 0.32 ;
        RECT  8.82 0.54 9.10 0.82 ;
        RECT  8.88 -0.28 9.04 0.82 ;
        RECT  7.78 0.54 8.06 0.82 ;
        RECT  7.84 -0.28 8.00 0.82 ;
        RECT  4.76 0.96 5.04 1.24 ;
        RECT  4.82 -0.28 4.98 1.24 ;
        RECT  0.10 0.96 0.38 1.24 ;
        RECT  0.16 -0.28 0.32 1.24 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.96 0.90 1.24 ;
        RECT  0.68 1.40 1.04 1.68 ;
        RECT  0.68 0.96 0.84 2.12 ;
        RECT  0.62 1.84 0.90 2.12 ;
        RECT  3.26 0.44 4.38 0.60 ;
        RECT  4.10 0.44 4.38 0.72 ;
        RECT  3.26 0.44 3.42 1.04 ;
        RECT  3.14 0.76 3.42 1.04 ;
        RECT  3.24 0.76 3.40 2.20 ;
        RECT  3.14 1.92 3.42 2.20 ;
        RECT  1.62 0.76 1.90 1.04 ;
        RECT  1.68 0.76 1.84 2.20 ;
        RECT  1.62 1.92 1.90 2.20 ;
        RECT  1.74 1.92 1.90 2.52 ;
        RECT  1.74 2.36 4.43 2.52 ;
        RECT  4.15 2.28 4.43 2.56 ;
        RECT  5.32 0.76 5.60 1.04 ;
        RECT  5.38 0.76 5.54 2.20 ;
        RECT  5.32 1.92 5.60 2.20 ;
        RECT  6.36 0.76 6.64 1.04 ;
        RECT  4.24 0.96 4.52 1.24 ;
        RECT  4.30 0.96 4.46 2.12 ;
        RECT  6.38 0.76 6.54 2.20 ;
        RECT  4.24 1.84 4.52 2.12 ;
        RECT  4.24 1.96 5.16 2.12 ;
        RECT  6.36 1.92 6.64 2.20 ;
        RECT  5.00 1.96 5.16 2.53 ;
        RECT  6.36 1.92 6.52 2.53 ;
        RECT  5.00 2.37 6.52 2.53 ;
        RECT  7.26 0.54 7.54 0.82 ;
        RECT  7.12 1.40 7.42 1.68 ;
        RECT  7.26 0.54 7.42 2.12 ;
        RECT  7.26 1.84 7.54 2.12 ;
        RECT  5.96 0.44 6.96 0.60 ;
        RECT  5.96 0.44 6.12 1.04 ;
        RECT  5.84 0.76 6.12 1.04 ;
        RECT  5.90 0.76 6.06 2.20 ;
        RECT  5.84 1.92 6.12 2.20 ;
        RECT  6.80 0.44 6.96 2.44 ;
        RECT  6.80 2.28 8.86 2.44 ;
        RECT  8.58 2.28 8.86 2.56 ;
    END
END MUX4LSP1V1_0

MACRO MUX3SP8V1_0
    CLASS CORE ;
    FOREIGN MUX3SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 13.23  LAYER ME1  ;
        ANTENNADIFFAREA 7.17  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.81  LAYER ME1  ;
        ANTENNAMAXAREACAR 16.41  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.98 1.84 7.26 2.12 ;
        RECT  6.98 0.96 7.26 1.24 ;
        RECT  6.98 0.96 7.14 2.12 ;
        RECT  6.14 1.52 7.14 1.68 ;
        RECT  6.14 0.96 6.30 1.98 ;
        RECT  5.94 2.26 6.22 2.54 ;
        RECT  6.06 1.82 6.22 2.54 ;
        RECT  5.94 0.96 6.30 1.24 ;
        END
    END OUT
    PIN B
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.18  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.58  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.12 1.92 2.42 2.20 ;
        RECT  2.12 0.76 2.42 1.04 ;
        RECT  2.06 1.46 2.34 1.74 ;
        RECT  2.12 0.76 2.28 2.20 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.52  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 22.68  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.20 1.46 1.54 1.74 ;
        RECT  1.10 1.92 1.38 2.20 ;
        RECT  1.10 0.76 1.38 1.04 ;
        RECT  1.20 0.76 1.36 2.20 ;
        END
    END A
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.90 1.40 3.32 1.68 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.33 0.44 1.75 ;
        END
    END S0
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.18 1.34 5.54 1.68 ;
        END
    END C
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 8.00 3.48 ;
        RECT  7.54 2.88 7.82 3.48 ;
        RECT  7.50 2.26 7.78 2.54 ;
        RECT  7.56 2.26 7.72 3.48 ;
        RECT  6.46 2.26 6.74 2.54 ;
        RECT  6.52 2.26 6.68 3.48 ;
        RECT  5.34 2.62 5.62 3.48 ;
        RECT  3.28 1.84 3.56 2.12 ;
        RECT  3.34 1.84 3.50 3.48 ;
        RECT  0.10 1.92 0.38 2.20 ;
        RECT  0.16 1.92 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 8.00 0.28 ;
        RECT  7.54 -0.28 7.82 0.32 ;
        RECT  7.50 0.54 7.78 0.82 ;
        RECT  7.56 -0.28 7.72 0.82 ;
        RECT  6.46 0.54 6.74 0.82 ;
        RECT  6.52 -0.28 6.68 0.82 ;
        RECT  5.42 0.68 5.70 0.96 ;
        RECT  5.48 -0.28 5.64 0.96 ;
        RECT  3.46 -0.28 3.74 0.68 ;
        RECT  0.10 0.76 0.38 1.04 ;
        RECT  0.16 -0.28 0.32 1.04 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.76 0.90 1.04 ;
        RECT  0.74 1.40 1.04 1.68 ;
        RECT  0.74 0.76 0.90 2.20 ;
        RECT  0.62 1.92 0.90 2.20 ;
        RECT  2.58 0.96 2.98 1.24 ;
        RECT  2.58 1.84 3.04 2.12 ;
        RECT  2.58 0.96 2.74 2.76 ;
        RECT  2.58 2.48 2.90 2.76 ;
        RECT  1.74 0.44 3.30 0.60 ;
        RECT  1.74 0.44 1.90 1.04 ;
        RECT  1.62 0.76 1.90 1.04 ;
        RECT  3.14 0.44 3.30 1.24 ;
        RECT  3.14 1.08 3.64 1.24 ;
        RECT  3.48 1.08 3.64 1.68 ;
        RECT  3.48 1.40 3.76 1.68 ;
        RECT  1.70 0.76 1.86 2.20 ;
        RECT  1.62 1.92 1.90 2.20 ;
        RECT  3.80 0.96 4.12 1.24 ;
        RECT  3.96 0.96 4.12 2.12 ;
        RECT  3.80 1.84 4.12 2.12 ;
        RECT  4.86 0.68 5.18 0.96 ;
        RECT  4.86 0.68 5.02 2.12 ;
        RECT  4.86 1.84 5.18 2.12 ;
        RECT  4.38 0.68 4.66 0.96 ;
        RECT  5.70 1.40 5.98 1.68 ;
        RECT  5.70 1.40 5.86 2.10 ;
        RECT  4.38 0.68 4.54 2.12 ;
        RECT  4.50 1.84 4.66 2.44 ;
        RECT  5.62 1.94 5.78 2.44 ;
        RECT  4.50 2.28 5.78 2.44 ;
    END
END MUX3SP8V1_0

MACRO MUX3SP4V1_0
    CLASS CORE ;
    FOREIGN MUX3SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.16 1.12 5.54 1.68 ;
        END
    END C
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.33 0.38 1.75 ;
        END
    END S0
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.90 1.40 3.24 1.70 ;
        END
    END S1
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.52  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 22.65  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.20 1.46 1.54 1.74 ;
        RECT  1.10 1.92 1.38 2.20 ;
        RECT  1.10 0.76 1.38 1.04 ;
        RECT  1.20 0.76 1.36 2.20 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.18  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.56  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.12 1.92 2.42 2.20 ;
        RECT  2.12 0.76 2.42 1.04 ;
        RECT  2.06 1.46 2.34 1.74 ;
        RECT  2.12 0.76 2.28 2.20 ;
        END
    END B
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 11.42  LAYER ME1  ;
        ANTENNADIFFAREA 5.49  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.42  LAYER ME1  ;
        ANTENNAMAXAREACAR 27.04  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.02 1.84 6.68 2.00 ;
        RECT  6.52 1.08 6.68 2.00 ;
        RECT  6.02 1.08 6.68 1.24 ;
        RECT  5.90 2.16 6.18 2.44 ;
        RECT  6.02 1.84 6.18 2.44 ;
        RECT  6.02 0.64 6.18 1.24 ;
        RECT  5.90 0.64 6.18 0.92 ;
        END
    END OUT
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 6.80 0.28 ;
        RECT  6.42 0.64 6.70 0.92 ;
        RECT  6.48 -0.28 6.64 0.92 ;
        RECT  6.34 -0.28 6.64 0.32 ;
        RECT  5.38 0.68 5.66 0.96 ;
        RECT  5.44 -0.28 5.60 0.96 ;
        RECT  3.42 -0.28 3.70 0.68 ;
        RECT  0.10 0.76 0.38 1.04 ;
        RECT  0.16 -0.28 0.32 1.04 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 6.80 3.48 ;
        RECT  6.42 2.16 6.70 2.44 ;
        RECT  6.34 2.88 6.64 3.48 ;
        RECT  6.48 2.16 6.64 3.48 ;
        RECT  5.30 2.62 5.58 3.48 ;
        RECT  3.18 1.86 3.46 2.14 ;
        RECT  3.24 1.86 3.40 3.48 ;
        RECT  0.10 1.92 0.38 2.20 ;
        RECT  0.16 1.92 0.32 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.76 0.90 1.04 ;
        RECT  0.74 1.40 1.04 1.68 ;
        RECT  0.74 0.76 0.90 2.20 ;
        RECT  0.62 1.92 0.90 2.20 ;
        RECT  2.58 0.96 2.94 1.24 ;
        RECT  2.58 1.86 2.94 2.14 ;
        RECT  2.58 0.96 2.74 2.76 ;
        RECT  2.52 2.48 2.80 2.76 ;
        RECT  1.74 0.44 3.26 0.60 ;
        RECT  1.74 0.44 1.90 1.04 ;
        RECT  1.62 0.76 1.90 1.04 ;
        RECT  3.10 0.44 3.26 1.24 ;
        RECT  3.10 1.08 3.56 1.24 ;
        RECT  3.40 1.08 3.56 1.68 ;
        RECT  3.40 1.40 3.72 1.68 ;
        RECT  1.70 0.76 1.86 2.20 ;
        RECT  1.62 1.92 1.90 2.20 ;
        RECT  3.72 0.96 4.04 1.24 ;
        RECT  3.88 0.96 4.04 2.14 ;
        RECT  3.74 1.86 4.04 2.14 ;
        RECT  4.84 0.68 5.14 0.96 ;
        RECT  4.84 0.68 5.00 2.14 ;
        RECT  4.84 1.86 5.14 2.14 ;
        RECT  4.30 0.68 4.62 0.96 ;
        RECT  5.70 1.40 5.98 1.68 ;
        RECT  5.70 1.40 5.86 2.00 ;
        RECT  4.30 0.68 4.46 2.14 ;
        RECT  4.46 1.86 4.62 2.44 ;
        RECT  5.58 1.84 5.74 2.44 ;
        RECT  4.46 2.28 5.74 2.44 ;
    END
END MUX3SP4V1_0

MACRO MUX3SP2V1_0
    CLASS CORE ;
    FOREIGN MUX3SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 10.53  LAYER ME1  ;
        ANTENNADIFFAREA 4.88  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.28  LAYER ME1  ;
        ANTENNAMAXAREACAR 37.82  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.00 1.84 6.32 2.12 ;
        RECT  6.16 0.96 6.32 2.12 ;
        RECT  6.00 0.96 6.32 1.24 ;
        END
    END OUT
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.24 1.12 5.52 1.68 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.19  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.67  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.14 1.92 2.42 2.20 ;
        RECT  2.14 0.76 2.42 1.04 ;
        RECT  2.06 1.46 2.34 1.74 ;
        RECT  2.14 0.76 2.30 2.20 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.52  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 22.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.22 1.46 1.54 1.74 ;
        RECT  1.10 1.92 1.38 2.20 ;
        RECT  1.22 0.76 1.38 2.20 ;
        RECT  1.10 0.76 1.38 1.04 ;
        END
    END A
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.90 1.40 3.32 1.68 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.40 0.50 1.68 ;
        END
    END S0
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 6.40 3.48 ;
        RECT  5.94 2.88 6.22 3.48 ;
        RECT  5.40 2.62 5.68 3.48 ;
        RECT  3.28 1.84 3.56 2.12 ;
        RECT  3.34 1.84 3.50 3.48 ;
        RECT  0.10 1.84 0.38 2.12 ;
        RECT  0.16 1.84 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 6.40 0.28 ;
        RECT  5.94 -0.28 6.22 0.32 ;
        RECT  5.48 0.68 5.76 0.96 ;
        RECT  5.54 -0.28 5.70 0.96 ;
        RECT  3.52 -0.28 3.80 0.68 ;
        RECT  0.10 0.96 0.38 1.24 ;
        RECT  0.16 -0.28 0.32 1.24 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.96 0.90 1.24 ;
        RECT  0.74 1.40 1.04 1.68 ;
        RECT  0.74 0.96 0.90 2.12 ;
        RECT  0.62 1.84 0.90 2.12 ;
        RECT  2.58 0.96 3.04 1.24 ;
        RECT  2.58 1.84 3.04 2.12 ;
        RECT  2.58 0.96 2.74 2.76 ;
        RECT  2.58 2.48 2.90 2.76 ;
        RECT  1.74 0.44 3.36 0.60 ;
        RECT  1.74 0.44 1.90 1.04 ;
        RECT  1.62 0.76 1.90 1.04 ;
        RECT  3.20 0.44 3.36 1.24 ;
        RECT  3.20 1.08 3.64 1.24 ;
        RECT  3.48 1.08 3.64 1.68 ;
        RECT  3.48 1.40 3.80 1.68 ;
        RECT  1.70 0.76 1.86 2.20 ;
        RECT  1.62 1.92 1.90 2.20 ;
        RECT  3.80 0.96 4.12 1.24 ;
        RECT  3.96 0.96 4.12 2.12 ;
        RECT  3.84 1.84 4.12 2.12 ;
        RECT  4.92 0.68 5.24 0.96 ;
        RECT  4.92 0.68 5.08 2.12 ;
        RECT  4.92 1.84 5.24 2.12 ;
        RECT  4.38 0.68 4.72 0.96 ;
        RECT  5.68 1.40 6.00 1.68 ;
        RECT  4.38 0.68 4.54 2.12 ;
        RECT  4.38 1.84 4.72 2.12 ;
        RECT  4.56 1.84 4.72 2.44 ;
        RECT  5.68 1.40 5.84 2.44 ;
        RECT  4.56 2.28 5.84 2.44 ;
    END
END MUX3SP2V1_0

MACRO MUX3SP1V1_0
    CLASS CORE ;
    FOREIGN MUX3SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.40 0.50 1.68 ;
        END
    END S0
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.90 1.40 3.32 1.68 ;
        END
    END S1
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.52  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 22.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.22 1.46 1.54 1.74 ;
        RECT  1.10 1.92 1.38 2.20 ;
        RECT  1.22 0.76 1.38 2.20 ;
        RECT  1.10 0.76 1.38 1.04 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.19  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.67  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.14 1.92 2.42 2.20 ;
        RECT  2.14 0.76 2.42 1.04 ;
        RECT  2.06 1.46 2.34 1.74 ;
        RECT  2.14 0.76 2.30 2.20 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.28 1.40 5.70 1.68 ;
        END
    END C
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 10.43  LAYER ME1  ;
        ANTENNADIFFAREA 4.52  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        ANTENNAMAXAREACAR 51.75  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.00 1.84 6.28 2.12 ;
        RECT  6.12 0.68 6.28 2.12 ;
        RECT  6.00 0.68 6.28 0.96 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 6.40 3.48 ;
        RECT  5.94 2.88 6.22 3.48 ;
        RECT  5.42 2.62 5.70 3.48 ;
        RECT  3.28 1.84 3.56 2.12 ;
        RECT  3.34 1.84 3.50 3.48 ;
        RECT  0.10 1.84 0.38 2.12 ;
        RECT  0.16 1.84 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 6.40 0.28 ;
        RECT  5.94 -0.28 6.22 0.32 ;
        RECT  5.48 0.68 5.76 0.96 ;
        RECT  5.54 -0.28 5.70 0.96 ;
        RECT  3.52 -0.28 3.80 0.68 ;
        RECT  0.10 0.96 0.38 1.24 ;
        RECT  0.16 -0.28 0.32 1.24 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.96 0.90 1.24 ;
        RECT  0.74 1.40 1.04 1.68 ;
        RECT  0.74 0.96 0.90 2.12 ;
        RECT  0.62 1.84 0.90 2.12 ;
        RECT  2.58 0.96 3.04 1.24 ;
        RECT  2.58 1.84 3.04 2.12 ;
        RECT  2.58 0.96 2.74 2.76 ;
        RECT  2.58 2.48 2.90 2.76 ;
        RECT  1.74 0.44 3.36 0.60 ;
        RECT  1.74 0.44 1.90 1.04 ;
        RECT  1.62 0.76 1.90 1.04 ;
        RECT  3.20 0.44 3.36 1.24 ;
        RECT  3.20 1.08 3.64 1.24 ;
        RECT  3.48 1.08 3.64 1.68 ;
        RECT  3.48 1.40 3.80 1.68 ;
        RECT  1.70 0.76 1.86 2.20 ;
        RECT  1.62 1.92 1.90 2.20 ;
        RECT  3.80 0.96 4.12 1.24 ;
        RECT  3.96 0.96 4.12 2.12 ;
        RECT  3.84 1.84 4.12 2.12 ;
        RECT  4.96 0.68 5.24 0.96 ;
        RECT  4.96 0.68 5.12 2.12 ;
        RECT  4.96 1.84 5.24 2.12 ;
        RECT  4.38 0.68 4.72 0.96 ;
        RECT  4.38 0.68 4.54 2.12 ;
        RECT  4.38 1.84 4.80 2.12 ;
        RECT  4.64 1.84 4.80 2.44 ;
        RECT  4.64 2.28 6.13 2.44 ;
        RECT  5.85 2.28 6.13 2.56 ;
    END
END MUX3SP1V1_0

MACRO MUX3ISP8V1_0
    CLASS CORE ;
    FOREIGN MUX3ISP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 22.31  LAYER ME1  ;
        ANTENNADIFFAREA 11.65  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.46  LAYER ME1  ;
        ANTENNAMAXAREACAR 15.29  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.78 1.84 12.06 2.12 ;
        RECT  8.66 1.08 12.06 1.24 ;
        RECT  11.78 0.96 12.06 1.24 ;
        RECT  10.74 1.84 12.06 2.00 ;
        RECT  11.32 1.08 11.48 2.00 ;
        RECT  10.74 1.84 11.02 2.12 ;
        RECT  10.74 0.96 11.02 1.24 ;
        RECT  9.70 0.96 9.98 1.24 ;
        RECT  8.66 0.96 8.94 1.24 ;
        END
    END OUT
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.44 1.26 2.72 1.68 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.90 1.34 2.28 1.68 ;
        END
    END S0
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.52 1.26 6.82 1.68 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.60  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 23.88  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.08 1.92 1.42 2.20 ;
        RECT  1.08 0.76 1.42 1.04 ;
        RECT  1.08 0.76 1.24 2.20 ;
        RECT  0.92 1.52 1.24 1.68 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.31  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 19.45  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.92 0.38 2.20 ;
        RECT  0.10 0.76 0.38 1.04 ;
        RECT  0.12 0.76 0.28 2.20 ;
        END
    END A
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 12.80 0.28 ;
        RECT  12.34 -0.28 12.62 0.32 ;
        RECT  12.30 0.62 12.58 0.90 ;
        RECT  12.36 -0.28 12.52 0.90 ;
        RECT  11.26 0.62 11.54 0.90 ;
        RECT  11.32 -0.28 11.48 0.90 ;
        RECT  10.22 0.62 10.50 0.90 ;
        RECT  10.28 -0.28 10.44 0.90 ;
        RECT  9.18 0.62 9.46 0.90 ;
        RECT  9.24 -0.28 9.40 0.90 ;
        RECT  8.14 0.62 8.42 0.90 ;
        RECT  8.20 -0.28 8.36 0.90 ;
        RECT  7.30 -0.28 7.58 0.58 ;
        RECT  5.20 0.96 5.48 1.24 ;
        RECT  5.26 -0.28 5.42 1.24 ;
        RECT  3.20 0.96 3.48 1.24 ;
        RECT  3.26 -0.28 3.42 1.24 ;
        RECT  2.14 0.82 2.42 1.10 ;
        RECT  2.20 -0.28 2.36 1.10 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 12.80 3.48 ;
        RECT  12.34 2.88 12.62 3.48 ;
        RECT  9.70 2.18 9.98 2.46 ;
        RECT  9.76 2.18 9.92 3.48 ;
        RECT  8.66 2.18 8.94 2.46 ;
        RECT  8.72 2.18 8.88 3.48 ;
        RECT  6.72 2.62 7.00 3.48 ;
        RECT  5.20 2.62 5.48 3.48 ;
        RECT  3.58 2.62 3.86 3.48 ;
        RECT  2.18 2.62 2.46 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  1.58 0.82 1.90 1.10 ;
        RECT  1.40 1.40 1.74 1.68 ;
        RECT  1.58 0.82 1.74 2.12 ;
        RECT  1.58 1.84 1.90 2.12 ;
        RECT  2.66 0.82 3.04 1.10 ;
        RECT  2.88 1.46 3.62 1.62 ;
        RECT  3.34 1.40 3.62 1.68 ;
        RECT  2.88 0.82 3.04 2.12 ;
        RECT  2.66 1.84 3.04 2.12 ;
        RECT  0.60 0.76 0.90 1.04 ;
        RECT  0.60 0.76 0.76 2.20 ;
        RECT  0.74 1.92 0.90 2.52 ;
        RECT  1.58 2.28 4.30 2.44 ;
        RECT  0.74 2.36 1.74 2.52 ;
        RECT  4.02 2.28 4.30 2.56 ;
        RECT  4.10 0.96 4.38 1.24 ;
        RECT  4.20 1.40 4.62 1.68 ;
        RECT  4.20 0.96 4.36 2.12 ;
        RECT  3.20 1.84 4.48 2.00 ;
        RECT  3.20 1.84 3.48 2.12 ;
        RECT  4.20 1.84 4.48 2.12 ;
        RECT  6.20 0.82 6.62 1.10 ;
        RECT  6.06 1.40 6.36 1.68 ;
        RECT  6.20 0.82 6.36 2.12 ;
        RECT  6.20 1.84 7.52 2.00 ;
        RECT  6.20 1.84 6.48 2.12 ;
        RECT  7.24 1.84 7.52 2.12 ;
        RECT  5.84 0.50 7.14 0.66 ;
        RECT  5.84 0.50 6.00 1.24 ;
        RECT  5.72 0.96 6.00 1.24 ;
        RECT  6.98 0.50 7.14 1.62 ;
        RECT  6.98 1.46 7.66 1.62 ;
        RECT  7.38 1.40 7.66 1.68 ;
        RECT  5.74 0.96 5.90 2.12 ;
        RECT  5.72 1.84 6.00 2.12 ;
        RECT  4.68 0.96 4.96 1.24 ;
        RECT  7.82 1.46 10.64 1.62 ;
        RECT  10.36 1.40 10.64 1.68 ;
        RECT  4.78 0.96 4.94 2.12 ;
        RECT  4.68 1.84 4.96 2.12 ;
        RECT  4.80 1.84 4.96 2.46 ;
        RECT  7.82 1.46 7.98 2.46 ;
        RECT  4.80 2.30 7.98 2.46 ;
        RECT  8.14 1.86 10.50 2.02 ;
        RECT  8.14 1.84 8.42 2.12 ;
        RECT  9.18 1.84 9.46 2.12 ;
        RECT  10.22 1.84 10.50 2.12 ;
        RECT  10.34 1.84 10.50 2.46 ;
        RECT  11.26 2.18 11.54 2.46 ;
        RECT  12.30 2.18 12.58 2.46 ;
        RECT  10.34 2.30 12.58 2.46 ;
    END
END MUX3ISP8V1_0

MACRO MUX3ISP4V1_0
    CLASS CORE ;
    FOREIGN MUX3ISP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 18.52  LAYER ME1  ;
        ANTENNADIFFAREA 9.10  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.88  LAYER ME1  ;
        ANTENNAMAXAREACAR 20.97  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.82 1.52 10.28 1.68 ;
        RECT  9.70 1.84 9.98 2.12 ;
        RECT  9.82 0.96 9.98 2.12 ;
        RECT  8.66 1.08 9.98 1.24 ;
        RECT  9.70 0.96 9.98 1.24 ;
        RECT  8.66 0.96 8.94 1.24 ;
        END
    END OUT
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.28  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 19.07  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.92 0.38 2.20 ;
        RECT  0.10 0.76 0.38 1.04 ;
        RECT  0.12 0.76 0.28 2.20 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.60  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 23.88  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.08 1.92 1.42 2.20 ;
        RECT  1.08 0.76 1.42 1.04 ;
        RECT  1.08 0.76 1.24 2.20 ;
        RECT  0.92 1.52 1.24 1.68 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.52 1.26 6.82 1.68 ;
        END
    END C
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.90 1.34 2.28 1.68 ;
        END
    END S0
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.44 1.26 2.72 1.68 ;
        END
    END S1
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 10.80 3.48 ;
        RECT  10.34 2.88 10.62 3.48 ;
        RECT  8.66 2.20 8.94 2.48 ;
        RECT  8.72 2.20 8.88 3.48 ;
        RECT  6.72 2.62 7.00 3.48 ;
        RECT  5.20 2.62 5.48 3.48 ;
        RECT  3.58 2.62 3.86 3.48 ;
        RECT  2.18 2.62 2.46 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 10.80 0.28 ;
        RECT  10.28 -0.28 10.62 0.32 ;
        RECT  10.22 0.60 10.50 0.88 ;
        RECT  10.28 -0.28 10.44 0.88 ;
        RECT  9.18 0.60 9.46 0.88 ;
        RECT  9.24 -0.28 9.40 0.88 ;
        RECT  8.14 0.60 8.42 0.88 ;
        RECT  8.20 -0.28 8.36 0.88 ;
        RECT  7.30 -0.28 7.58 0.58 ;
        RECT  5.20 0.96 5.48 1.24 ;
        RECT  5.26 -0.28 5.42 1.24 ;
        RECT  3.20 0.96 3.48 1.24 ;
        RECT  3.26 -0.28 3.42 1.24 ;
        RECT  2.14 0.82 2.42 1.10 ;
        RECT  2.20 -0.28 2.36 1.10 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  1.58 0.82 1.90 1.10 ;
        RECT  1.40 1.40 1.74 1.68 ;
        RECT  1.58 0.82 1.74 2.12 ;
        RECT  1.58 1.84 1.90 2.12 ;
        RECT  2.66 0.82 3.04 1.10 ;
        RECT  2.88 1.46 3.62 1.62 ;
        RECT  3.34 1.40 3.62 1.68 ;
        RECT  2.88 0.82 3.04 2.12 ;
        RECT  2.66 1.84 3.04 2.12 ;
        RECT  0.60 0.76 0.90 1.04 ;
        RECT  0.60 0.76 0.76 2.20 ;
        RECT  0.74 1.92 0.90 2.52 ;
        RECT  1.58 2.28 4.30 2.44 ;
        RECT  0.74 2.36 1.74 2.52 ;
        RECT  4.02 2.28 4.30 2.56 ;
        RECT  4.10 0.96 4.38 1.24 ;
        RECT  4.20 1.40 4.62 1.68 ;
        RECT  4.20 0.96 4.36 2.12 ;
        RECT  3.20 1.84 4.48 2.00 ;
        RECT  3.20 1.84 3.48 2.12 ;
        RECT  4.20 1.84 4.48 2.12 ;
        RECT  6.20 0.82 6.62 1.10 ;
        RECT  6.06 1.40 6.36 1.68 ;
        RECT  6.20 0.82 6.36 2.12 ;
        RECT  6.20 1.84 7.52 2.00 ;
        RECT  6.20 1.84 6.48 2.12 ;
        RECT  7.24 1.84 7.52 2.12 ;
        RECT  5.84 0.50 7.14 0.66 ;
        RECT  5.84 0.50 6.00 1.24 ;
        RECT  5.72 0.96 6.00 1.24 ;
        RECT  6.98 0.50 7.14 1.62 ;
        RECT  6.98 1.46 7.66 1.62 ;
        RECT  7.38 1.40 7.66 1.68 ;
        RECT  5.74 0.96 5.90 2.12 ;
        RECT  5.72 1.84 6.00 2.12 ;
        RECT  4.68 0.96 4.96 1.24 ;
        RECT  7.82 1.46 9.60 1.62 ;
        RECT  9.32 1.40 9.60 1.68 ;
        RECT  4.78 0.96 4.94 2.12 ;
        RECT  4.68 1.84 4.96 2.12 ;
        RECT  4.80 1.84 4.96 2.46 ;
        RECT  7.82 1.46 7.98 2.46 ;
        RECT  4.80 2.30 7.98 2.46 ;
        RECT  8.14 1.88 9.46 2.04 ;
        RECT  8.14 1.84 8.42 2.12 ;
        RECT  9.18 1.84 9.46 2.12 ;
        RECT  9.30 1.84 9.46 2.48 ;
        RECT  10.22 2.20 10.50 2.48 ;
        RECT  9.30 2.32 10.50 2.48 ;
    END
END MUX3ISP4V1_0

MACRO MUX3ISP2V1_0
    CLASS CORE ;
    FOREIGN MUX3ISP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 16.04  LAYER ME1  ;
        ANTENNADIFFAREA 7.33  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER ME1  ;
        ANTENNAMAXAREACAR 28.33  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.78 1.08 9.10 1.24 ;
        RECT  8.82 0.96 9.10 1.24 ;
        RECT  7.85 1.84 8.27 2.12 ;
        RECT  8.11 1.08 8.27 2.12 ;
        RECT  7.78 0.96 8.06 1.24 ;
        RECT  7.78 0.66 7.94 1.24 ;
        RECT  7.68 0.66 7.94 0.94 ;
        END
    END OUT
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.44 1.26 2.72 1.68 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.90 1.34 2.28 1.68 ;
        END
    END S0
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.48 1.26 6.76 1.68 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.68  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 25.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.06 1.92 1.42 2.20 ;
        RECT  1.06 0.76 1.42 1.04 ;
        RECT  1.06 0.76 1.22 2.20 ;
        RECT  0.86 1.46 1.22 1.74 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.38  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 20.57  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.92 0.38 2.20 ;
        RECT  0.10 0.76 0.38 1.04 ;
        RECT  0.12 0.76 0.28 2.20 ;
        END
    END A
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 9.20 0.28 ;
        RECT  8.74 -0.28 9.02 0.32 ;
        RECT  8.30 0.62 8.58 0.90 ;
        RECT  8.36 -0.28 8.52 0.90 ;
        RECT  7.24 0.82 7.52 1.10 ;
        RECT  7.30 -0.28 7.46 1.10 ;
        RECT  5.20 0.96 5.48 1.24 ;
        RECT  5.26 -0.28 5.42 1.24 ;
        RECT  3.20 0.96 3.48 1.24 ;
        RECT  3.26 -0.28 3.42 1.24 ;
        RECT  2.14 0.82 2.42 1.10 ;
        RECT  2.20 -0.28 2.36 1.10 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 9.20 3.48 ;
        RECT  8.75 2.18 9.03 2.46 ;
        RECT  8.74 2.88 9.02 3.48 ;
        RECT  8.81 2.18 8.97 3.48 ;
        RECT  6.72 2.62 7.00 3.48 ;
        RECT  5.20 2.62 5.48 3.48 ;
        RECT  3.58 2.62 3.86 3.48 ;
        RECT  2.18 2.62 2.46 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  1.58 0.82 1.90 1.10 ;
        RECT  1.40 1.40 1.74 1.68 ;
        RECT  1.58 0.82 1.74 2.12 ;
        RECT  1.58 1.84 1.90 2.12 ;
        RECT  2.66 0.82 3.04 1.10 ;
        RECT  2.88 1.46 3.62 1.62 ;
        RECT  3.34 1.40 3.62 1.68 ;
        RECT  2.88 0.82 3.04 2.12 ;
        RECT  2.66 1.84 3.04 2.12 ;
        RECT  0.54 0.76 0.90 1.04 ;
        RECT  0.54 0.76 0.70 2.20 ;
        RECT  0.54 1.92 0.90 2.20 ;
        RECT  0.74 1.92 0.90 2.52 ;
        RECT  1.58 2.28 4.30 2.44 ;
        RECT  0.74 2.36 1.74 2.52 ;
        RECT  4.02 2.28 4.30 2.56 ;
        RECT  4.10 0.96 4.38 1.24 ;
        RECT  4.20 1.40 4.62 1.68 ;
        RECT  4.20 0.96 4.36 2.12 ;
        RECT  3.20 1.84 4.48 2.00 ;
        RECT  3.20 1.84 3.48 2.12 ;
        RECT  4.20 1.84 4.48 2.12 ;
        RECT  6.16 0.82 6.62 1.10 ;
        RECT  6.00 1.40 6.32 1.68 ;
        RECT  6.16 0.82 6.32 2.12 ;
        RECT  6.16 1.84 7.52 2.00 ;
        RECT  6.16 1.84 6.48 2.12 ;
        RECT  7.24 1.84 7.52 2.12 ;
        RECT  5.84 0.50 7.08 0.66 ;
        RECT  5.84 0.50 6.00 1.24 ;
        RECT  6.92 0.50 7.08 1.62 ;
        RECT  6.92 1.46 7.91 1.62 ;
        RECT  7.63 1.40 7.91 1.68 ;
        RECT  5.68 0.96 5.84 2.12 ;
        RECT  5.68 1.84 6.00 2.12 ;
        RECT  4.68 0.96 4.96 1.24 ;
        RECT  8.51 1.40 8.79 1.68 ;
        RECT  4.78 0.96 4.94 2.12 ;
        RECT  4.68 1.84 4.96 2.12 ;
        RECT  4.80 1.84 4.96 2.46 ;
        RECT  8.43 1.45 8.59 2.46 ;
        RECT  4.80 2.30 8.59 2.46 ;
    END
END MUX3ISP2V1_0

MACRO MUX3ISP1V1_0
    CLASS CORE ;
    FOREIGN MUX3ISP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.28  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 19.07  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.92 0.38 2.20 ;
        RECT  0.10 0.76 0.38 1.04 ;
        RECT  0.12 0.76 0.28 2.20 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.60  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 23.88  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.08 1.92 1.42 2.20 ;
        RECT  1.08 0.76 1.42 1.04 ;
        RECT  1.08 0.76 1.24 2.20 ;
        RECT  0.92 1.52 1.24 1.68 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.52 1.26 6.82 1.68 ;
        END
    END C
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.90 1.34 2.28 1.68 ;
        END
    END S0
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.44 1.26 2.72 1.68 ;
        END
    END S1
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 15.65  LAYER ME1  ;
        ANTENNADIFFAREA 7.05  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.40  LAYER ME1  ;
        ANTENNAMAXAREACAR 38.82  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.69 1.84 9.08 2.12 ;
        RECT  8.92 0.96 9.08 2.12 ;
        RECT  8.76 0.96 9.08 1.24 ;
        RECT  7.72 1.02 9.08 1.18 ;
        RECT  7.72 0.96 8.00 1.24 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 9.20 3.48 ;
        RECT  8.74 2.88 9.02 3.48 ;
        RECT  7.64 2.62 7.92 3.48 ;
        RECT  6.72 2.62 7.00 3.48 ;
        RECT  5.20 2.62 5.48 3.48 ;
        RECT  3.58 2.62 3.86 3.48 ;
        RECT  2.18 2.62 2.46 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 9.20 0.28 ;
        RECT  8.74 -0.28 9.02 0.32 ;
        RECT  8.24 -0.28 8.52 0.58 ;
        RECT  7.30 -0.28 7.58 0.58 ;
        RECT  5.20 0.96 5.48 1.24 ;
        RECT  5.26 -0.28 5.42 1.24 ;
        RECT  3.20 0.96 3.48 1.24 ;
        RECT  3.26 -0.28 3.42 1.24 ;
        RECT  2.14 0.82 2.42 1.10 ;
        RECT  2.20 -0.28 2.36 1.10 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  1.58 0.82 1.90 1.10 ;
        RECT  1.40 1.40 1.74 1.68 ;
        RECT  1.58 0.82 1.74 2.12 ;
        RECT  1.58 1.84 1.90 2.12 ;
        RECT  2.66 0.82 3.04 1.10 ;
        RECT  2.88 1.46 3.62 1.62 ;
        RECT  3.34 1.40 3.62 1.68 ;
        RECT  2.88 0.82 3.04 2.12 ;
        RECT  2.66 1.84 3.04 2.12 ;
        RECT  0.60 0.76 0.90 1.04 ;
        RECT  0.60 0.76 0.76 2.20 ;
        RECT  0.74 1.92 0.90 2.52 ;
        RECT  1.58 2.28 4.30 2.44 ;
        RECT  0.74 2.36 1.74 2.52 ;
        RECT  4.02 2.28 4.30 2.56 ;
        RECT  4.10 0.96 4.38 1.24 ;
        RECT  4.20 1.40 4.62 1.68 ;
        RECT  4.20 0.96 4.36 2.12 ;
        RECT  3.20 1.84 4.48 2.00 ;
        RECT  3.20 1.84 3.48 2.12 ;
        RECT  4.20 1.84 4.48 2.12 ;
        RECT  6.20 0.82 6.62 1.10 ;
        RECT  6.06 1.40 6.36 1.68 ;
        RECT  6.20 0.82 6.36 2.12 ;
        RECT  6.20 1.84 7.52 2.00 ;
        RECT  6.20 1.84 6.48 2.12 ;
        RECT  7.24 1.84 7.52 2.12 ;
        RECT  4.68 0.96 4.96 1.24 ;
        RECT  4.78 0.96 4.94 2.12 ;
        RECT  4.68 1.84 4.96 2.12 ;
        RECT  4.80 1.84 4.96 2.46 ;
        RECT  4.80 2.30 8.31 2.46 ;
        RECT  8.03 2.22 8.31 2.50 ;
        RECT  5.84 0.50 7.14 0.66 ;
        RECT  5.84 0.50 6.00 1.24 ;
        RECT  5.72 0.96 6.00 1.24 ;
        RECT  6.98 0.50 7.14 1.62 ;
        RECT  6.98 1.46 8.73 1.62 ;
        RECT  8.45 1.40 8.73 1.68 ;
        RECT  5.74 0.96 5.90 2.12 ;
        RECT  5.72 1.84 6.00 2.12 ;
    END
END MUX3ISP1V1_0

MACRO MUX2SP8V1_0
    CLASS CORE ;
    FOREIGN MUX2SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.42 1.26 2.70 1.68 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.90 1.26 1.18 1.68 ;
        END
    END B
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.42 1.26 0.70 1.68 ;
        END
    END S
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 9.51  LAYER ME1  ;
        ANTENNADIFFAREA 5.62  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER ME1  ;
        ANTENNAMAXAREACAR 13.96  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.28 1.84 4.56 2.12 ;
        RECT  4.28 0.96 4.56 1.24 ;
        RECT  4.28 0.96 4.44 2.12 ;
        RECT  3.34 1.52 4.44 1.68 ;
        RECT  3.24 1.84 3.52 2.12 ;
        RECT  3.24 0.96 3.52 1.24 ;
        RECT  3.34 0.96 3.50 2.12 ;
        END
    END OUT
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 5.20 0.28 ;
        RECT  4.80 0.64 5.08 0.92 ;
        RECT  4.86 -0.28 5.02 0.92 ;
        RECT  4.74 -0.28 5.02 0.32 ;
        RECT  3.76 0.64 4.04 0.92 ;
        RECT  3.82 -0.28 3.98 0.92 ;
        RECT  2.72 0.68 3.00 0.96 ;
        RECT  2.78 -0.28 2.94 0.96 ;
        RECT  0.62 0.68 0.90 0.96 ;
        RECT  0.68 -0.28 0.84 0.96 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 5.20 3.48 ;
        RECT  4.80 2.16 5.08 2.44 ;
        RECT  4.74 2.88 5.02 3.48 ;
        RECT  4.86 2.16 5.02 3.48 ;
        RECT  3.76 2.16 4.04 2.44 ;
        RECT  3.82 2.16 3.98 3.48 ;
        RECT  2.66 2.62 2.94 3.48 ;
        RECT  0.40 2.52 0.68 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  1.14 0.68 1.50 0.96 ;
        RECT  1.34 0.68 1.50 2.12 ;
        RECT  1.14 1.84 1.50 2.12 ;
        RECT  0.10 0.68 0.38 0.96 ;
        RECT  0.10 0.68 0.26 2.12 ;
        RECT  0.10 1.90 0.98 2.06 ;
        RECT  0.10 1.84 0.38 2.12 ;
        RECT  0.82 1.90 0.98 2.44 ;
        RECT  0.82 2.28 1.60 2.44 ;
        RECT  1.32 2.28 1.60 2.56 ;
        RECT  2.10 0.68 2.48 0.96 ;
        RECT  2.10 0.68 2.26 2.12 ;
        RECT  2.10 1.84 2.48 2.12 ;
        RECT  1.66 0.68 1.94 0.96 ;
        RECT  2.90 1.40 3.18 1.68 ;
        RECT  1.72 0.68 1.88 2.12 ;
        RECT  1.66 1.84 1.94 2.12 ;
        RECT  1.78 1.84 1.94 2.44 ;
        RECT  2.90 1.40 3.06 2.44 ;
        RECT  1.78 2.28 3.06 2.44 ;
    END
END MUX2SP8V1_0

MACRO MUX2SP4V1_0
    CLASS CORE ;
    FOREIGN MUX2SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 7.70  LAYER ME1  ;
        ANTENNADIFFAREA 4.26  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.36  LAYER ME1  ;
        ANTENNAMAXAREACAR 21.69  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.34 1.52 3.88 1.68 ;
        RECT  3.24 1.84 3.52 2.12 ;
        RECT  3.24 0.96 3.52 1.24 ;
        RECT  3.34 0.96 3.50 2.12 ;
        END
    END OUT
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.42 1.26 0.70 1.68 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.90 1.26 1.18 1.68 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.42 1.26 2.70 1.68 ;
        END
    END A
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.40 3.48 ;
        RECT  3.82 2.88 4.22 3.48 ;
        RECT  3.76 2.16 4.04 2.44 ;
        RECT  3.82 2.16 3.98 3.48 ;
        RECT  2.66 2.62 2.94 3.48 ;
        RECT  0.40 2.52 0.68 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.40 0.28 ;
        RECT  3.82 -0.28 4.22 0.32 ;
        RECT  3.76 0.64 4.04 0.92 ;
        RECT  3.82 -0.28 3.98 0.92 ;
        RECT  2.72 0.68 3.00 0.96 ;
        RECT  2.78 -0.28 2.94 0.96 ;
        RECT  0.62 0.68 0.90 0.96 ;
        RECT  0.68 -0.28 0.84 0.96 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  1.14 0.68 1.50 0.96 ;
        RECT  1.34 0.68 1.50 2.12 ;
        RECT  1.14 1.84 1.50 2.12 ;
        RECT  0.10 0.68 0.38 0.96 ;
        RECT  0.10 0.68 0.26 2.12 ;
        RECT  0.10 1.90 0.98 2.06 ;
        RECT  0.10 1.84 0.38 2.12 ;
        RECT  0.82 1.90 0.98 2.44 ;
        RECT  0.82 2.28 1.60 2.44 ;
        RECT  1.32 2.28 1.60 2.56 ;
        RECT  2.10 0.68 2.48 0.96 ;
        RECT  2.10 0.68 2.26 2.12 ;
        RECT  2.10 1.84 2.48 2.12 ;
        RECT  1.66 0.68 1.94 0.96 ;
        RECT  2.90 1.40 3.18 1.68 ;
        RECT  1.72 0.68 1.88 2.12 ;
        RECT  1.66 1.84 1.94 2.12 ;
        RECT  1.78 1.84 1.94 2.44 ;
        RECT  2.90 1.40 3.06 2.44 ;
        RECT  1.78 2.28 3.06 2.44 ;
    END
END MUX2SP4V1_0

MACRO MUX2SP2V1_0
    CLASS CORE ;
    FOREIGN MUX2SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.42 1.26 2.70 1.68 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.90 1.26 1.18 1.68 ;
        END
    END B
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.42 1.26 0.70 1.68 ;
        END
    END S
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 7.34  LAYER ME1  ;
        ANTENNADIFFAREA 3.66  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.21  LAYER ME1  ;
        ANTENNAMAXAREACAR 34.73  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.36 1.46 3.92 1.74 ;
        RECT  3.24 1.84 3.52 2.12 ;
        RECT  3.36 0.96 3.52 2.12 ;
        RECT  3.24 0.96 3.52 1.24 ;
        END
    END OUT
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.00 0.28 ;
        RECT  3.54 -0.28 3.82 0.32 ;
        RECT  2.72 0.68 3.00 0.96 ;
        RECT  2.78 -0.28 2.94 0.96 ;
        RECT  0.62 0.68 0.90 0.96 ;
        RECT  0.68 -0.28 0.84 0.96 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.00 3.48 ;
        RECT  3.54 2.88 3.82 3.48 ;
        RECT  2.64 2.62 2.92 3.48 ;
        RECT  0.40 2.52 0.68 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  1.14 0.68 1.50 0.96 ;
        RECT  1.34 0.68 1.50 2.12 ;
        RECT  1.14 1.84 1.50 2.12 ;
        RECT  0.10 0.68 0.38 0.96 ;
        RECT  0.10 0.68 0.26 2.12 ;
        RECT  0.10 1.90 0.98 2.06 ;
        RECT  0.10 1.84 0.38 2.12 ;
        RECT  0.82 1.90 0.98 2.44 ;
        RECT  0.82 2.28 1.60 2.44 ;
        RECT  1.32 2.28 1.60 2.56 ;
        RECT  2.10 0.68 2.48 0.96 ;
        RECT  2.10 0.68 2.26 2.12 ;
        RECT  2.10 1.84 2.48 2.12 ;
        RECT  1.66 0.68 1.94 0.96 ;
        RECT  2.88 1.40 3.18 1.68 ;
        RECT  1.72 0.68 1.88 2.12 ;
        RECT  1.66 1.84 1.94 2.12 ;
        RECT  1.78 1.84 1.94 2.44 ;
        RECT  2.88 1.40 3.04 2.44 ;
        RECT  1.78 2.28 3.04 2.44 ;
    END
END MUX2SP2V1_0

MACRO MUX2SP1V1_0
    CLASS CORE ;
    FOREIGN MUX2SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.48 1.26 2.76 1.68 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.90 1.26 1.18 1.68 ;
        END
    END B
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.42 1.26 0.70 1.68 ;
        END
    END S
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 6.39  LAYER ME1  ;
        ANTENNADIFFAREA 3.13  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        ANTENNAMAXAREACAR 47.51  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.22 1.84 3.50 2.12 ;
        RECT  3.22 0.68 3.50 0.96 ;
        RECT  3.32 0.68 3.48 2.12 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 3.60 3.48 ;
        RECT  3.14 2.88 3.42 3.48 ;
        RECT  2.64 2.61 2.92 3.48 ;
        RECT  0.40 2.52 0.68 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 3.60 0.28 ;
        RECT  3.14 -0.28 3.42 0.32 ;
        RECT  2.70 0.68 2.98 0.96 ;
        RECT  2.76 -0.28 2.92 0.96 ;
        RECT  0.62 0.68 0.90 0.96 ;
        RECT  0.68 -0.28 0.84 0.96 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  1.14 0.68 1.50 0.96 ;
        RECT  1.34 0.68 1.50 2.12 ;
        RECT  1.14 1.84 1.50 2.12 ;
        RECT  0.10 0.68 0.38 0.96 ;
        RECT  0.10 0.68 0.26 2.12 ;
        RECT  0.10 1.90 0.98 2.06 ;
        RECT  0.10 1.84 0.38 2.12 ;
        RECT  0.82 1.90 0.98 2.44 ;
        RECT  0.82 2.28 1.60 2.44 ;
        RECT  1.32 2.28 1.60 2.56 ;
        RECT  2.16 0.68 2.46 0.96 ;
        RECT  2.16 0.68 2.32 2.12 ;
        RECT  2.16 1.84 2.46 2.12 ;
        RECT  1.66 0.68 1.94 0.96 ;
        RECT  1.72 0.68 1.88 2.12 ;
        RECT  1.66 1.84 1.94 2.12 ;
        RECT  1.78 1.84 1.94 2.44 ;
        RECT  1.78 2.28 3.36 2.44 ;
        RECT  3.08 2.28 3.36 2.56 ;
    END
END MUX2SP1V1_0

MACRO MUX2LSP8V1_0
    CLASS CORE ;
    FOREIGN MUX2LSP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 15.40  LAYER ME1  ;
        ANTENNADIFFAREA 9.41  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.76  LAYER ME1  ;
        ANTENNAMAXAREACAR 20.30  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.37 1.84 7.65 2.12 ;
        RECT  4.25 1.08 7.65 1.24 ;
        RECT  7.37 0.96 7.65 1.24 ;
        RECT  6.33 1.84 7.65 2.00 ;
        RECT  6.46 1.08 6.74 2.00 ;
        RECT  6.33 1.84 6.61 2.12 ;
        RECT  6.33 0.96 6.61 1.24 ;
        RECT  5.29 0.96 5.57 1.24 ;
        RECT  4.25 0.96 4.53 1.24 ;
        END
    END OUT
    PIN EN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.69  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.60 1.40 8.02 1.68 ;
        END
    END EN
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.46 1.34 0.74 1.76 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.76 1.06 3.18 1.34 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.90 1.46 1.32 1.76 ;
        END
    END A
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 8.80 0.28 ;
        RECT  8.34 -0.28 8.62 0.32 ;
        RECT  7.89 0.52 8.17 0.80 ;
        RECT  7.95 -0.28 8.11 0.80 ;
        RECT  6.85 0.52 7.13 0.80 ;
        RECT  6.91 -0.28 7.07 0.80 ;
        RECT  5.81 0.52 6.09 0.80 ;
        RECT  5.87 -0.28 6.03 0.80 ;
        RECT  4.77 0.52 5.05 0.80 ;
        RECT  4.83 -0.28 4.99 0.80 ;
        RECT  3.73 0.52 4.01 0.80 ;
        RECT  3.79 -0.28 3.95 0.80 ;
        RECT  2.98 0.62 3.26 0.90 ;
        RECT  3.04 -0.28 3.20 0.90 ;
        RECT  0.86 0.76 1.14 1.04 ;
        RECT  0.92 -0.28 1.08 1.04 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 8.80 3.48 ;
        RECT  8.34 2.88 8.62 3.48 ;
        RECT  5.29 2.28 5.57 2.56 ;
        RECT  5.35 2.28 5.51 3.48 ;
        RECT  4.25 2.28 4.53 2.56 ;
        RECT  4.31 2.28 4.47 3.48 ;
        RECT  3.39 2.62 3.67 3.48 ;
        RECT  0.86 1.92 1.14 2.20 ;
        RECT  0.92 1.92 1.08 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.14 0.76 0.62 1.04 ;
        RECT  0.14 0.76 0.30 2.20 ;
        RECT  0.14 1.92 0.62 2.20 ;
        RECT  0.26 1.92 0.42 2.76 ;
        RECT  0.20 2.48 0.48 2.76 ;
        RECT  1.38 0.76 1.66 1.04 ;
        RECT  1.50 0.76 1.66 2.20 ;
        RECT  1.38 1.92 1.66 2.20 ;
        RECT  2.44 0.62 2.74 0.90 ;
        RECT  2.44 0.62 2.60 2.20 ;
        RECT  2.44 1.92 2.74 2.20 ;
        RECT  1.90 0.76 2.18 1.04 ;
        RECT  4.07 1.40 4.35 1.68 ;
        RECT  3.08 1.52 4.35 1.68 ;
        RECT  1.96 0.76 2.12 2.20 ;
        RECT  1.90 1.92 2.18 2.20 ;
        RECT  2.02 1.92 2.18 2.52 ;
        RECT  3.08 1.52 3.24 2.52 ;
        RECT  2.02 2.36 3.24 2.52 ;
        RECT  3.73 1.90 6.09 2.06 ;
        RECT  3.73 1.84 4.01 2.12 ;
        RECT  4.77 1.84 5.05 2.12 ;
        RECT  5.81 1.84 6.09 2.12 ;
        RECT  5.93 1.84 6.09 2.56 ;
        RECT  6.85 2.28 7.13 2.56 ;
        RECT  7.89 2.28 8.17 2.56 ;
        RECT  5.93 2.40 8.17 2.56 ;
    END
END MUX2LSP8V1_0

MACRO MUX2LSP4V1_0
    CLASS CORE ;
    FOREIGN MUX2LSP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.90 1.46 1.32 1.74 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.76 1.08 3.18 1.36 ;
        END
    END B
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.46 1.34 0.74 1.76 ;
        END
    END S
    PIN EN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.31  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.79 1.40 5.21 1.68 ;
        END
    END EN
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 11.41  LAYER ME1  ;
        ANTENNADIFFAREA 6.07  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.38  LAYER ME1  ;
        ANTENNAMAXAREACAR 30.29  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.40 1.46 5.94 1.74 ;
        RECT  5.28 1.84 5.56 2.12 ;
        RECT  5.40 0.91 5.56 2.12 ;
        RECT  4.24 1.03 5.56 1.19 ;
        RECT  5.28 0.91 5.56 1.19 ;
        RECT  4.24 0.91 4.52 1.19 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 6.40 3.48 ;
        RECT  5.94 2.88 6.22 3.48 ;
        RECT  4.24 2.20 4.52 2.48 ;
        RECT  4.30 2.20 4.46 3.48 ;
        RECT  3.43 2.62 3.71 3.48 ;
        RECT  0.86 1.92 1.14 2.20 ;
        RECT  0.92 1.92 1.08 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 6.40 0.28 ;
        RECT  5.86 -0.28 6.22 0.32 ;
        RECT  5.80 0.54 6.08 0.82 ;
        RECT  5.86 -0.28 6.02 0.82 ;
        RECT  4.76 0.54 5.04 0.82 ;
        RECT  4.82 -0.28 4.98 0.82 ;
        RECT  3.72 0.54 4.00 0.82 ;
        RECT  3.78 -0.28 3.94 0.82 ;
        RECT  2.98 0.64 3.26 0.92 ;
        RECT  3.04 -0.28 3.20 0.92 ;
        RECT  0.86 0.76 1.14 1.04 ;
        RECT  0.92 -0.28 1.08 1.04 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.14 0.76 0.62 1.04 ;
        RECT  0.14 0.76 0.30 2.20 ;
        RECT  0.14 1.92 0.62 2.20 ;
        RECT  0.26 1.92 0.42 2.76 ;
        RECT  0.20 2.48 0.48 2.76 ;
        RECT  1.38 0.76 1.66 1.04 ;
        RECT  1.50 0.76 1.66 2.20 ;
        RECT  1.38 1.92 1.66 2.20 ;
        RECT  2.44 0.64 2.74 0.92 ;
        RECT  2.44 0.64 2.60 2.20 ;
        RECT  2.44 1.92 2.74 2.20 ;
        RECT  1.90 0.76 2.18 1.04 ;
        RECT  4.24 1.40 4.52 1.68 ;
        RECT  3.14 1.52 4.52 1.68 ;
        RECT  1.96 0.76 2.12 2.20 ;
        RECT  1.90 1.92 2.18 2.20 ;
        RECT  2.02 1.92 2.18 2.52 ;
        RECT  3.14 1.52 3.30 2.52 ;
        RECT  2.02 2.36 3.30 2.52 ;
        RECT  3.72 1.84 4.92 2.00 ;
        RECT  3.72 1.84 4.00 2.12 ;
        RECT  4.76 1.84 4.92 2.46 ;
        RECT  4.76 2.18 5.04 2.46 ;
        RECT  5.80 2.18 6.08 2.46 ;
        RECT  4.76 2.30 6.08 2.46 ;
    END
END MUX2LSP4V1_0

MACRO MUX2LSP2V1_0
    CLASS CORE ;
    FOREIGN MUX2LSP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 8.51  LAYER ME1  ;
        ANTENNADIFFAREA 4.35  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.22  LAYER ME1  ;
        ANTENNAMAXAREACAR 39.41  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.02 1.84 4.68 2.12 ;
        RECT  4.52 1.00 4.68 2.12 ;
        RECT  3.50 1.00 4.68 1.16 ;
        RECT  3.50 0.88 3.78 1.16 ;
        END
    END OUT
    PIN EN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.15  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.26 1.40 3.54 1.82 ;
        END
    END EN
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.46 1.34 0.74 1.76 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.66 1.40 3.10 1.68 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.90 1.46 1.32 1.76 ;
        END
    END A
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.80 0.28 ;
        RECT  4.08 -0.28 4.62 0.32 ;
        RECT  4.02 0.54 4.30 0.82 ;
        RECT  4.08 -0.28 4.24 0.82 ;
        RECT  2.94 -0.28 3.22 0.58 ;
        RECT  0.86 0.76 1.14 1.04 ;
        RECT  0.92 -0.28 1.08 1.04 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.80 3.48 ;
        RECT  4.34 2.88 4.62 3.48 ;
        RECT  2.89 2.62 3.17 3.48 ;
        RECT  0.86 1.92 1.14 2.20 ;
        RECT  0.92 1.92 1.08 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.14 0.76 0.62 1.04 ;
        RECT  0.14 0.76 0.30 2.20 ;
        RECT  0.14 1.92 0.62 2.20 ;
        RECT  0.26 1.92 0.42 2.76 ;
        RECT  0.20 2.48 0.48 2.76 ;
        RECT  1.38 0.76 1.66 1.04 ;
        RECT  1.50 0.76 1.66 2.20 ;
        RECT  1.38 1.92 1.66 2.20 ;
        RECT  2.34 0.88 2.74 1.16 ;
        RECT  2.34 0.86 2.50 2.12 ;
        RECT  2.34 1.84 2.74 2.12 ;
        RECT  1.90 0.76 2.18 1.04 ;
        RECT  3.70 1.40 4.02 1.68 ;
        RECT  1.96 0.76 2.12 2.20 ;
        RECT  1.90 1.92 2.18 2.20 ;
        RECT  2.02 1.92 2.18 2.44 ;
        RECT  3.70 1.40 3.86 2.44 ;
        RECT  2.02 2.28 3.86 2.44 ;
    END
END MUX2LSP2V1_0

MACRO MUX2LSP1V1_0
    CLASS CORE ;
    FOREIGN MUX2LSP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.92 1.48 1.34 1.76 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.66 1.40 3.08 1.68 ;
        END
    END B
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.48 1.34 0.76 1.76 ;
        END
    END S
    PIN EN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.26 1.12 3.54 1.54 ;
        END
    END EN
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 7.85  LAYER ME1  ;
        ANTENNADIFFAREA 3.46  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        ANTENNAMAXAREACAR 58.38  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.88 1.84 4.16 2.12 ;
        RECT  3.88 1.52 4.04 2.12 ;
        RECT  3.70 1.52 4.04 1.68 ;
        RECT  3.70 0.68 3.86 1.68 ;
        RECT  3.50 0.68 3.86 0.96 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.40 3.48 ;
        RECT  3.94 2.88 4.22 3.48 ;
        RECT  2.89 2.62 3.17 3.48 ;
        RECT  0.86 1.92 1.14 2.20 ;
        RECT  0.92 1.92 1.08 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.40 0.28 ;
        RECT  4.02 0.68 4.30 0.96 ;
        RECT  4.08 -0.28 4.24 0.96 ;
        RECT  3.94 -0.28 4.24 0.32 ;
        RECT  2.98 0.68 3.26 0.96 ;
        RECT  3.04 -0.28 3.20 0.96 ;
        RECT  0.86 0.76 1.14 1.04 ;
        RECT  0.92 -0.28 1.08 1.04 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.16 0.76 0.62 1.04 ;
        RECT  0.16 0.76 0.32 2.20 ;
        RECT  0.16 1.92 0.62 2.20 ;
        RECT  0.26 1.92 0.42 2.76 ;
        RECT  0.20 2.48 0.48 2.76 ;
        RECT  1.38 0.76 1.66 1.04 ;
        RECT  1.50 0.76 1.66 2.20 ;
        RECT  1.38 1.92 1.66 2.20 ;
        RECT  2.34 0.68 2.74 0.96 ;
        RECT  2.34 0.68 2.50 2.12 ;
        RECT  2.34 1.84 2.74 2.12 ;
        RECT  1.90 0.76 2.18 1.04 ;
        RECT  1.96 0.76 2.12 2.20 ;
        RECT  1.90 1.92 2.18 2.20 ;
        RECT  2.02 1.92 2.18 2.44 ;
        RECT  2.02 2.28 3.94 2.44 ;
        RECT  3.66 2.28 3.94 2.56 ;
    END
END MUX2LSP1V1_0

MACRO MUX2ISP8V1_0
    CLASS CORE ;
    FOREIGN MUX2ISP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 9.01  LAYER ME1  ;
        ANTENNADIFFAREA 4.80  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 134.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.26 1.84 4.54 2.48 ;
        RECT  4.26 0.60 4.54 1.24 ;
        RECT  4.26 0.60 4.42 2.48 ;
        RECT  3.32 1.52 4.42 1.68 ;
        RECT  3.22 1.84 3.50 2.48 ;
        RECT  3.22 0.60 3.50 1.24 ;
        RECT  3.32 0.60 3.48 2.48 ;
        END
    END OUT
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.40 0.50 1.68 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.12  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.61  LAYER ME1  ;
        ANTENNAMAXAREACAR 1.83  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.14 1.92 2.42 2.20 ;
        RECT  2.14 0.76 2.42 1.04 ;
        RECT  2.20 0.76 2.36 2.20 ;
        RECT  2.12 1.52 2.36 1.68 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.14  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.61  LAYER ME1  ;
        ANTENNAMAXAREACAR 1.86  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.20 1.52 1.48 1.68 ;
        RECT  1.10 1.92 1.38 2.20 ;
        RECT  1.10 0.76 1.38 1.04 ;
        RECT  1.20 0.76 1.36 2.20 ;
        END
    END A
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 5.20 3.48 ;
        RECT  4.78 1.84 5.06 2.48 ;
        RECT  4.74 2.88 5.02 3.48 ;
        RECT  4.84 1.84 5.00 3.48 ;
        RECT  3.74 1.84 4.02 2.48 ;
        RECT  3.80 1.84 3.96 3.48 ;
        RECT  2.70 1.84 2.98 2.48 ;
        RECT  2.76 1.84 2.92 3.48 ;
        RECT  0.10 1.84 0.38 2.12 ;
        RECT  0.16 1.84 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 5.20 0.28 ;
        RECT  4.78 0.60 5.06 1.24 ;
        RECT  4.74 -0.28 5.02 0.32 ;
        RECT  4.84 -0.28 5.00 1.24 ;
        RECT  3.74 0.60 4.02 1.24 ;
        RECT  3.80 -0.28 3.96 1.24 ;
        RECT  2.70 0.60 2.98 1.24 ;
        RECT  2.76 -0.28 2.92 1.24 ;
        RECT  0.10 0.96 0.38 1.24 ;
        RECT  0.16 -0.28 0.32 1.24 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.96 0.90 1.24 ;
        RECT  0.68 1.40 1.04 1.68 ;
        RECT  0.68 0.96 0.84 2.12 ;
        RECT  0.62 1.84 0.90 2.12 ;
        RECT  1.62 0.76 1.90 1.04 ;
        RECT  1.62 1.92 1.90 2.20 ;
        RECT  1.68 0.76 1.84 2.64 ;
        RECT  1.68 2.48 2.54 2.64 ;
        RECT  2.26 2.48 2.54 2.76 ;
    END
END MUX2ISP8V1_0

MACRO MUX2ISP4V1_0
    CLASS CORE ;
    FOREIGN MUX2ISP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 7.07  LAYER ME1  ;
        ANTENNADIFFAREA 3.31  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 105.14  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.22 1.84 3.50 2.48 ;
        RECT  3.22 0.60 3.50 1.24 ;
        RECT  3.32 0.60 3.48 2.48 ;
        END
    END OUT
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.13  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.31  LAYER ME1  ;
        ANTENNAMAXAREACAR 3.67  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.20 1.52 1.48 1.68 ;
        RECT  1.10 1.92 1.38 2.20 ;
        RECT  1.10 0.76 1.38 1.04 ;
        RECT  1.20 0.76 1.36 2.20 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.83  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.31  LAYER ME1  ;
        ANTENNAMAXAREACAR 2.70  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.14 1.92 2.42 2.20 ;
        RECT  2.14 0.76 2.42 1.04 ;
        RECT  2.20 0.76 2.36 2.20 ;
        RECT  2.12 1.52 2.36 1.68 ;
        END
    END B
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.40 0.50 1.68 ;
        END
    END S
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.40 0.28 ;
        RECT  3.80 -0.28 4.22 0.32 ;
        RECT  3.74 0.60 4.02 1.24 ;
        RECT  3.80 -0.28 3.96 1.24 ;
        RECT  2.70 0.60 2.98 1.24 ;
        RECT  2.76 -0.28 2.92 1.24 ;
        RECT  0.10 0.96 0.38 1.24 ;
        RECT  0.16 -0.28 0.32 1.24 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.40 3.48 ;
        RECT  3.80 2.88 4.22 3.48 ;
        RECT  3.74 1.84 4.02 2.48 ;
        RECT  3.80 1.84 3.96 3.48 ;
        RECT  2.70 1.84 2.98 2.48 ;
        RECT  2.76 1.84 2.92 3.48 ;
        RECT  0.10 1.84 0.38 2.12 ;
        RECT  0.16 1.84 0.32 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.96 0.90 1.24 ;
        RECT  0.68 1.40 1.04 1.68 ;
        RECT  0.68 0.96 0.84 2.12 ;
        RECT  0.62 1.84 0.90 2.12 ;
        RECT  1.62 0.76 1.90 1.04 ;
        RECT  1.62 1.92 1.90 2.20 ;
        RECT  1.68 0.76 1.84 2.64 ;
        RECT  1.68 2.48 2.54 2.64 ;
        RECT  2.26 2.48 2.54 2.76 ;
    END
END MUX2ISP4V1_0

MACRO MUX2ISP2V1_0
    CLASS CORE ;
    FOREIGN MUX2ISP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 5.69  LAYER ME1  ;
        ANTENNADIFFAREA 2.51  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 84.65  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.76 1.52 3.08 1.68 ;
        RECT  2.70 1.84 2.98 2.46 ;
        RECT  2.70 0.62 2.98 1.24 ;
        RECT  2.76 0.62 2.92 2.46 ;
        END
    END OUT
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.40 0.50 1.68 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.12  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.15  LAYER ME1  ;
        ANTENNAMAXAREACAR 7.54  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.14 1.92 2.42 2.20 ;
        RECT  2.14 0.76 2.42 1.04 ;
        RECT  2.20 0.76 2.36 2.20 ;
        RECT  2.12 1.52 2.36 1.68 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.14  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.15  LAYER ME1  ;
        ANTENNAMAXAREACAR 7.67  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.20 1.52 1.48 1.68 ;
        RECT  1.10 1.92 1.38 2.20 ;
        RECT  1.10 0.76 1.38 1.04 ;
        RECT  1.20 0.76 1.36 2.20 ;
        END
    END A
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 3.60 0.28 ;
        RECT  3.22 0.62 3.50 1.24 ;
        RECT  3.27 -0.28 3.43 1.24 ;
        RECT  3.14 -0.28 3.43 0.32 ;
        RECT  0.10 0.96 0.38 1.24 ;
        RECT  0.16 -0.28 0.32 1.24 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 3.60 3.48 ;
        RECT  3.22 1.84 3.50 2.46 ;
        RECT  3.14 2.88 3.42 3.48 ;
        RECT  3.26 1.84 3.42 3.48 ;
        RECT  0.10 1.84 0.38 2.12 ;
        RECT  0.16 1.84 0.32 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.96 0.90 1.24 ;
        RECT  0.68 1.40 1.04 1.68 ;
        RECT  0.68 0.96 0.84 2.12 ;
        RECT  0.62 1.84 0.90 2.12 ;
        RECT  1.62 0.76 1.90 1.04 ;
        RECT  1.62 1.92 1.90 2.20 ;
        RECT  1.68 0.76 1.84 2.64 ;
        RECT  1.68 2.48 2.54 2.64 ;
        RECT  2.26 2.48 2.54 2.76 ;
    END
END MUX2ISP2V1_0

MACRO MUX2ISP1V1_0
    CLASS CORE ;
    FOREIGN MUX2ISP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.19  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.69  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.20 1.52 1.48 1.68 ;
        RECT  1.10 1.92 1.38 2.20 ;
        RECT  1.10 0.76 1.38 1.04 ;
        RECT  1.20 0.76 1.36 2.20 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.89  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 13.26  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.14 1.92 2.42 2.20 ;
        RECT  2.14 0.76 2.42 1.04 ;
        RECT  2.20 0.76 2.36 2.20 ;
        RECT  2.12 1.52 2.36 1.68 ;
        END
    END B
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.40 0.50 1.68 ;
        END
    END S
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 5.14  LAYER ME1  ;
        ANTENNADIFFAREA 2.05  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 76.45  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.64 1.84 2.92 2.12 ;
        RECT  2.64 0.96 2.92 1.24 ;
        RECT  2.68 0.96 2.84 2.12 ;
        RECT  2.52 1.52 2.84 1.68 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 3.60 3.48 ;
        RECT  3.16 1.84 3.44 2.12 ;
        RECT  3.14 2.88 3.42 3.48 ;
        RECT  3.26 1.84 3.42 3.48 ;
        RECT  0.10 1.84 0.38 2.12 ;
        RECT  0.16 1.84 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 3.60 0.28 ;
        RECT  3.16 0.96 3.44 1.24 ;
        RECT  3.14 -0.28 3.42 0.32 ;
        RECT  3.22 -0.28 3.38 1.24 ;
        RECT  0.10 0.96 0.38 1.24 ;
        RECT  0.16 -0.28 0.32 1.24 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.96 0.90 1.24 ;
        RECT  0.68 1.40 1.04 1.68 ;
        RECT  0.68 0.96 0.84 2.12 ;
        RECT  0.62 1.84 0.90 2.12 ;
        RECT  1.62 0.76 1.90 1.04 ;
        RECT  1.68 0.76 1.84 2.20 ;
        RECT  1.62 1.92 1.90 2.20 ;
        RECT  1.74 1.92 1.90 2.52 ;
        RECT  1.74 2.36 3.10 2.52 ;
        RECT  2.82 2.28 3.10 2.56 ;
    END
END MUX2ISP1V1_0

MACRO MA2OF3SP8V1_0
    CLASS CORE ;
    FOREIGN MA2OF3SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 9.89  LAYER ME1  ;
        ANTENNADIFFAREA 5.93  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.58  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.18  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.14 1.98 4.42 2.58 ;
        RECT  4.14 0.62 4.42 1.22 ;
        RECT  4.14 0.62 4.30 2.58 ;
        RECT  3.22 1.52 4.30 1.68 ;
        RECT  3.22 1.46 3.54 1.74 ;
        RECT  3.10 1.98 3.38 2.58 ;
        RECT  3.22 0.62 3.38 2.58 ;
        RECT  3.10 0.62 3.38 1.22 ;
        END
    END OUT
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.46 1.46 1.94 1.74 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.80 1.44 1.20 1.76 ;
        END
    END IN3
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.44 0.44 1.76 ;
        END
    END IN1
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 5.20 0.28 ;
        RECT  4.72 -0.28 5.02 0.32 ;
        RECT  4.66 0.62 4.94 1.22 ;
        RECT  4.72 -0.28 4.88 1.22 ;
        RECT  3.62 0.62 3.90 1.22 ;
        RECT  3.68 -0.28 3.84 1.22 ;
        RECT  2.58 0.62 2.86 1.22 ;
        RECT  2.64 -0.28 2.80 1.22 ;
        RECT  0.62 0.68 0.90 0.96 ;
        RECT  0.68 -0.28 0.84 0.96 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 5.20 3.48 ;
        RECT  4.72 2.88 5.02 3.48 ;
        RECT  4.66 1.98 4.94 2.58 ;
        RECT  4.72 1.98 4.88 3.48 ;
        RECT  3.62 1.98 3.90 2.58 ;
        RECT  3.68 1.98 3.84 3.48 ;
        RECT  2.58 1.98 2.86 2.58 ;
        RECT  2.64 1.98 2.80 3.48 ;
        RECT  0.62 2.24 0.90 2.52 ;
        RECT  0.68 2.24 0.84 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.21 1.92 1.30 2.08 ;
        RECT  0.21 1.92 0.37 2.52 ;
        RECT  1.14 1.92 1.30 2.52 ;
        RECT  0.10 2.24 0.38 2.52 ;
        RECT  1.14 2.24 1.42 2.52 ;
        RECT  0.10 0.68 0.38 0.96 ;
        RECT  1.14 0.68 1.42 0.96 ;
        RECT  0.22 0.68 0.38 1.28 ;
        RECT  1.14 0.68 1.30 1.28 ;
        RECT  0.22 1.12 1.30 1.28 ;
        RECT  1.66 0.68 1.94 0.96 ;
        RECT  1.78 0.68 1.94 1.28 ;
        RECT  1.78 1.12 2.26 1.28 ;
        RECT  2.10 1.52 3.02 1.68 ;
        RECT  2.74 1.46 3.02 1.74 ;
        RECT  2.10 1.12 2.26 2.08 ;
        RECT  1.78 1.92 2.26 2.08 ;
        RECT  1.78 1.92 1.94 2.52 ;
        RECT  1.66 2.24 1.94 2.52 ;
    END
END MA2OF3SP8V1_0

MACRO MA2OF3SP4V1_0
    CLASS CORE ;
    FOREIGN MA2OF3SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.44 0.44 1.76 ;
        END
    END IN1
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.80 1.44 1.20 1.76 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.46 1.46 1.94 1.74 ;
        END
    END IN2
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 7.55  LAYER ME1  ;
        ANTENNADIFFAREA 4.11  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.29  LAYER ME1  ;
        ANTENNAMAXAREACAR 26.22  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.22 1.46 3.54 1.74 ;
        RECT  3.10 1.98 3.38 2.58 ;
        RECT  3.22 0.62 3.38 2.58 ;
        RECT  3.10 0.62 3.38 1.22 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.00 3.48 ;
        RECT  3.62 1.98 3.90 2.58 ;
        RECT  3.54 2.88 3.84 3.48 ;
        RECT  3.68 1.98 3.84 3.48 ;
        RECT  2.58 1.98 2.86 2.58 ;
        RECT  2.64 1.98 2.80 3.48 ;
        RECT  0.62 2.24 0.90 2.52 ;
        RECT  0.68 2.24 0.84 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.00 0.28 ;
        RECT  3.62 0.62 3.90 1.22 ;
        RECT  3.68 -0.28 3.84 1.22 ;
        RECT  3.54 -0.28 3.84 0.32 ;
        RECT  2.58 0.62 2.86 1.22 ;
        RECT  2.64 -0.28 2.80 1.22 ;
        RECT  0.62 0.68 0.90 0.96 ;
        RECT  0.68 -0.28 0.84 0.96 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.21 1.92 1.30 2.08 ;
        RECT  0.21 1.92 0.37 2.52 ;
        RECT  1.14 1.92 1.30 2.52 ;
        RECT  0.10 2.24 0.38 2.52 ;
        RECT  1.14 2.24 1.42 2.52 ;
        RECT  0.10 0.68 0.38 0.96 ;
        RECT  1.14 0.68 1.42 0.96 ;
        RECT  0.22 0.68 0.38 1.28 ;
        RECT  1.14 0.68 1.30 1.28 ;
        RECT  0.22 1.12 1.30 1.28 ;
        RECT  1.66 0.68 1.94 0.96 ;
        RECT  1.78 0.68 1.94 1.28 ;
        RECT  1.78 1.12 2.26 1.28 ;
        RECT  2.10 1.52 3.02 1.68 ;
        RECT  2.74 1.46 3.02 1.74 ;
        RECT  2.10 1.12 2.26 2.08 ;
        RECT  1.78 1.92 2.26 2.08 ;
        RECT  1.78 1.92 1.94 2.52 ;
        RECT  1.66 2.24 1.94 2.52 ;
    END
END MA2OF3SP4V1_0

MACRO MA2OF3SP2V1_0
    CLASS CORE ;
    FOREIGN MA2OF3SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 6.72  LAYER ME1  ;
        ANTENNADIFFAREA 3.28  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.14  LAYER ME1  ;
        ANTENNAMAXAREACAR 46.67  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.12 1.98 3.48 2.58 ;
        RECT  3.32 0.62 3.48 2.58 ;
        RECT  3.12 0.62 3.48 1.22 ;
        END
    END OUT
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.46 1.46 1.94 1.74 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.80 1.44 1.20 1.76 ;
        END
    END IN3
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.44 0.44 1.76 ;
        END
    END IN1
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 3.60 0.28 ;
        RECT  3.14 -0.28 3.42 0.32 ;
        RECT  2.60 0.62 2.88 1.22 ;
        RECT  2.66 -0.28 2.82 1.22 ;
        RECT  0.62 0.68 0.90 0.96 ;
        RECT  0.68 -0.28 0.84 0.96 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 3.60 3.48 ;
        RECT  3.14 2.88 3.42 3.48 ;
        RECT  2.60 1.98 2.88 2.58 ;
        RECT  2.66 1.98 2.82 3.48 ;
        RECT  0.62 2.24 0.90 2.52 ;
        RECT  0.68 2.24 0.84 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.21 1.92 1.30 2.08 ;
        RECT  0.21 1.92 0.37 2.52 ;
        RECT  1.14 1.92 1.30 2.52 ;
        RECT  0.10 2.24 0.38 2.52 ;
        RECT  1.14 2.24 1.42 2.52 ;
        RECT  0.10 0.68 0.38 0.96 ;
        RECT  1.14 0.68 1.42 0.96 ;
        RECT  0.22 0.68 0.38 1.28 ;
        RECT  1.14 0.68 1.30 1.28 ;
        RECT  0.22 1.12 1.30 1.28 ;
        RECT  1.66 0.68 1.94 0.96 ;
        RECT  1.78 0.68 1.94 1.28 ;
        RECT  1.78 1.12 2.26 1.28 ;
        RECT  2.10 1.52 3.02 1.68 ;
        RECT  2.74 1.46 3.02 1.74 ;
        RECT  2.10 1.12 2.26 2.08 ;
        RECT  1.78 1.92 2.26 2.08 ;
        RECT  1.78 1.92 1.94 2.52 ;
        RECT  1.66 2.24 1.94 2.52 ;
    END
END MA2OF3SP2V1_0

MACRO MA2OF3SP1V1_0
    CLASS CORE ;
    FOREIGN MA2OF3SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 6.52  LAYER ME1  ;
        ANTENNADIFFAREA 2.82  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 96.99  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.08 2.24 3.48 2.52 ;
        RECT  3.32 0.68 3.48 2.52 ;
        RECT  3.08 0.68 3.48 0.96 ;
        END
    END OUT
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.46 1.46 1.94 1.74 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.44 0.44 1.76 ;
        END
    END IN1
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.80 1.44 1.20 1.76 ;
        END
    END IN3
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 3.60 3.48 ;
        RECT  3.14 2.88 3.42 3.48 ;
        RECT  2.56 2.24 2.84 2.52 ;
        RECT  2.62 2.24 2.78 3.48 ;
        RECT  0.62 2.24 0.90 2.52 ;
        RECT  0.68 2.24 0.84 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 3.60 0.28 ;
        RECT  3.14 -0.28 3.42 0.32 ;
        RECT  2.56 0.68 2.84 0.96 ;
        RECT  2.62 -0.28 2.78 0.96 ;
        RECT  0.62 0.68 0.90 0.96 ;
        RECT  0.68 -0.28 0.84 0.96 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.21 1.92 1.30 2.08 ;
        RECT  0.21 1.92 0.37 2.52 ;
        RECT  1.14 1.92 1.30 2.52 ;
        RECT  0.10 2.24 0.38 2.52 ;
        RECT  1.14 2.24 1.42 2.52 ;
        RECT  0.10 0.68 0.38 0.96 ;
        RECT  1.14 0.68 1.42 0.96 ;
        RECT  0.22 0.68 0.38 1.28 ;
        RECT  1.14 0.68 1.30 1.28 ;
        RECT  0.22 1.12 1.30 1.28 ;
        RECT  1.66 0.68 1.94 0.96 ;
        RECT  1.78 0.68 1.94 1.28 ;
        RECT  1.78 1.12 2.88 1.28 ;
        RECT  2.72 1.46 3.02 1.74 ;
        RECT  2.72 1.12 2.88 2.08 ;
        RECT  1.78 1.92 2.88 2.08 ;
        RECT  1.78 1.92 1.94 2.52 ;
        RECT  1.66 2.24 1.94 2.52 ;
    END
END MA2OF3SP1V1_0

MACRO INVTSP8V1_0
    CLASS CORE ;
    FOREIGN INVTSP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 10.63  LAYER ME1  ;
        ANTENNADIFFAREA 7.22  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.34  LAYER ME1  ;
        ANTENNAMAXAREACAR 31.65  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.92 1.90 5.20 2.18 ;
        RECT  4.92 0.96 5.20 1.24 ;
        RECT  4.92 0.96 5.08 2.18 ;
        RECT  4.00 1.52 5.08 1.68 ;
        RECT  3.88 1.90 4.16 2.18 ;
        RECT  4.00 0.96 4.16 2.18 ;
        RECT  3.88 0.96 4.16 1.24 ;
        END
    END OUT
    PIN IN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.54  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.14 1.46 1.54 1.74 ;
        END
    END IN
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.45  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.42 1.46 0.84 1.74 ;
        END
    END E
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 6.00 3.48 ;
        RECT  5.54 2.88 5.82 3.48 ;
        RECT  2.88 2.22 3.16 2.50 ;
        RECT  2.94 2.22 3.10 3.48 ;
        RECT  1.84 2.22 2.12 2.50 ;
        RECT  1.90 2.22 2.06 3.48 ;
        RECT  0.80 2.22 1.08 2.50 ;
        RECT  0.86 2.22 1.02 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 6.00 0.28 ;
        RECT  5.54 -0.28 5.82 0.32 ;
        RECT  2.88 0.68 3.16 0.96 ;
        RECT  2.94 -0.28 3.10 0.96 ;
        RECT  1.84 0.68 2.12 0.96 ;
        RECT  1.90 -0.28 2.06 0.96 ;
        RECT  0.80 0.68 1.08 0.96 ;
        RECT  0.86 -0.28 1.02 0.96 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.96 0.52 1.24 ;
        RECT  0.10 0.96 0.26 2.76 ;
        RECT  0.10 2.10 0.52 2.38 ;
        RECT  0.10 2.10 0.38 2.76 ;
        RECT  1.32 1.90 3.64 2.06 ;
        RECT  3.36 1.90 3.64 2.18 ;
        RECT  1.32 1.90 1.60 2.22 ;
        RECT  2.36 1.90 2.64 2.22 ;
        RECT  3.48 1.90 3.64 2.50 ;
        RECT  3.48 2.34 5.72 2.50 ;
        RECT  4.40 2.32 4.68 2.60 ;
        RECT  5.44 2.32 5.72 2.60 ;
        RECT  3.48 0.64 5.72 0.80 ;
        RECT  4.40 0.54 4.68 0.82 ;
        RECT  5.44 0.54 5.72 0.82 ;
        RECT  1.32 0.96 1.60 1.28 ;
        RECT  2.36 0.96 2.64 1.28 ;
        RECT  3.36 0.96 3.64 1.28 ;
        RECT  3.48 0.64 3.64 1.28 ;
        RECT  1.32 1.12 3.64 1.28 ;
    END
END INVTSP8V1_0

MACRO INVTSP4V1_0
    CLASS CORE ;
    FOREIGN INVTSP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.28  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.42 1.46 0.84 1.74 ;
        END
    END E
    PIN IN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.27  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.14 1.46 1.54 1.74 ;
        END
    END IN
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 6.64  LAYER ME1  ;
        ANTENNADIFFAREA 4.57  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.17  LAYER ME1  ;
        ANTENNAMAXAREACAR 39.51  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.84 1.90 3.12 2.18 ;
        RECT  2.84 0.96 3.12 1.24 ;
        RECT  2.92 0.96 3.08 2.18 ;
        END
    END OUT
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.00 0.28 ;
        RECT  3.54 -0.28 3.82 0.32 ;
        RECT  1.84 0.68 2.12 0.96 ;
        RECT  1.90 -0.28 2.06 0.96 ;
        RECT  0.80 0.68 1.08 0.96 ;
        RECT  0.86 -0.28 1.02 0.96 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.00 3.48 ;
        RECT  3.54 2.88 3.82 3.48 ;
        RECT  1.84 2.22 2.12 2.50 ;
        RECT  1.90 2.22 2.06 3.48 ;
        RECT  0.80 2.22 1.08 2.50 ;
        RECT  0.86 2.22 1.02 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.96 0.52 1.24 ;
        RECT  0.10 0.96 0.26 2.76 ;
        RECT  0.10 2.10 0.52 2.38 ;
        RECT  0.10 2.10 0.38 2.76 ;
        RECT  1.32 1.90 2.60 2.06 ;
        RECT  2.32 1.90 2.60 2.18 ;
        RECT  1.32 1.90 1.60 2.22 ;
        RECT  2.44 1.90 2.60 2.50 ;
        RECT  2.44 2.34 3.64 2.50 ;
        RECT  3.36 2.32 3.64 2.60 ;
        RECT  2.44 0.64 3.64 0.80 ;
        RECT  3.36 0.54 3.64 0.82 ;
        RECT  1.32 0.96 1.60 1.28 ;
        RECT  2.32 0.96 2.60 1.28 ;
        RECT  2.44 0.64 2.60 1.28 ;
        RECT  1.32 1.12 2.60 1.28 ;
    END
END INVTSP4V1_0

MACRO INVTSP2V1_0
    CLASS CORE ;
    FOREIGN INVTSP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 2.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 3.51  LAYER ME1  ;
        ANTENNADIFFAREA 2.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.08  LAYER ME1  ;
        ANTENNAMAXAREACAR 41.78  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.72 1.96 2.08 2.24 ;
        RECT  1.72 0.96 2.08 1.24 ;
        RECT  1.72 0.96 1.88 2.24 ;
        END
    END OUT
    PIN IN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.12  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.10 1.46 1.54 1.74 ;
        END
    END IN
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.42 1.46 0.84 1.74 ;
        END
    END E
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 2.40 3.48 ;
        RECT  1.94 2.88 2.22 3.48 ;
        RECT  0.76 2.10 1.04 2.38 ;
        RECT  0.82 2.10 0.98 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 2.40 0.28 ;
        RECT  1.94 -0.28 2.22 0.32 ;
        RECT  0.76 0.76 1.04 1.04 ;
        RECT  0.82 -0.28 0.98 1.04 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.96 0.52 1.24 ;
        RECT  0.10 0.96 0.26 2.76 ;
        RECT  0.10 2.10 0.52 2.38 ;
        RECT  0.10 2.10 0.38 2.76 ;
    END
END INVTSP2V1_0

MACRO INVTSP1V1_0
    CLASS CORE ;
    FOREIGN INVTSP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 2.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 3.15  LAYER ME1  ;
        ANTENNADIFFAREA 1.49  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.03  LAYER ME1  ;
        ANTENNAMAXAREACAR 93.76  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.46 2.36 1.88 2.64 ;
        RECT  1.72 0.56 1.88 2.64 ;
        RECT  1.46 0.56 1.88 0.84 ;
        END
    END OUT
    PIN IN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.80 1.48 1.22 1.76 ;
        END
    END IN
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.10  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.28 1.04 1.56 1.32 ;
        RECT  0.44 1.12 1.56 1.28 ;
        RECT  0.44 1.06 0.72 1.34 ;
        END
    END E
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 2.00 3.48 ;
        RECT  1.54 2.88 1.82 3.48 ;
        RECT  0.62 2.36 0.90 2.64 ;
        RECT  0.68 2.36 0.84 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 2.00 0.28 ;
        RECT  1.54 -0.28 1.82 0.32 ;
        RECT  0.62 0.56 0.90 0.84 ;
        RECT  0.68 -0.28 0.84 0.84 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.56 0.38 0.84 ;
        RECT  0.10 1.92 1.56 2.08 ;
        RECT  1.28 1.92 1.56 2.20 ;
        RECT  0.10 0.56 0.26 2.64 ;
        RECT  0.10 2.36 0.38 2.64 ;
    END
END INVTSP1V1_0

MACRO INVSP8V1_0
    CLASS CORE ;
    FOREIGN INVSP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 2.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 4.54  LAYER ME1  ;
        ANTENNADIFFAREA 3.29  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.66 1.90 1.94 2.50 ;
        RECT  1.66 0.64 1.94 1.24 ;
        RECT  1.66 0.64 1.82 2.50 ;
        RECT  0.74 1.52 1.82 1.68 ;
        RECT  0.74 1.46 1.14 1.74 ;
        RECT  0.62 1.90 0.90 2.50 ;
        RECT  0.74 0.64 0.90 2.50 ;
        RECT  0.62 0.64 0.90 1.24 ;
        END
    END OUT
    PIN IN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.58  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.46 0.56 1.74 ;
        END
    END IN
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 2.80 3.48 ;
        RECT  2.24 2.88 2.62 3.48 ;
        RECT  2.18 1.90 2.46 2.50 ;
        RECT  2.24 1.90 2.40 3.48 ;
        RECT  1.14 1.90 1.42 2.50 ;
        RECT  1.20 1.90 1.36 3.48 ;
        RECT  0.10 1.90 0.38 2.50 ;
        RECT  0.16 1.90 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 2.80 0.28 ;
        RECT  2.24 -0.28 2.62 0.32 ;
        RECT  2.18 0.64 2.46 1.24 ;
        RECT  2.24 -0.28 2.40 1.24 ;
        RECT  1.14 0.64 1.42 1.24 ;
        RECT  1.20 -0.28 1.36 1.24 ;
        RECT  0.10 0.64 0.38 1.24 ;
        RECT  0.16 -0.28 0.32 1.24 ;
        END
    END GND!
END INVSP8V1_0

MACRO INVSP6V1_0
    CLASS CORE ;
    FOREIGN INVSP6V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 2.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.43  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.46 0.64 1.74 ;
        END
    END IN
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 3.63  LAYER ME1  ;
        ANTENNADIFFAREA 2.68  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.74 1.90 2.02 2.50 ;
        RECT  1.74 0.64 2.02 1.24 ;
        RECT  1.74 0.64 1.90 2.50 ;
        RECT  0.82 1.52 1.90 1.68 ;
        RECT  0.82 1.46 1.14 1.74 ;
        RECT  0.70 1.90 0.98 2.50 ;
        RECT  0.82 0.64 0.98 2.50 ;
        RECT  0.70 0.64 0.98 1.24 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 2.40 3.48 ;
        RECT  1.94 2.88 2.22 3.48 ;
        RECT  1.22 1.90 1.50 2.50 ;
        RECT  1.28 1.90 1.44 3.48 ;
        RECT  0.18 1.90 0.46 2.50 ;
        RECT  0.24 1.90 0.40 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 2.40 0.28 ;
        RECT  1.94 -0.28 2.22 0.32 ;
        RECT  1.22 0.64 1.50 1.24 ;
        RECT  1.28 -0.28 1.44 1.24 ;
        RECT  0.18 0.64 0.46 1.24 ;
        RECT  0.24 -0.28 0.40 1.24 ;
        END
    END GND!
END INVSP6V1_0

MACRO INVSP64V1_0
    CLASS CORE ;
    FOREIGN INVSP64V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 17.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 4.61  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.46 0.56 1.74 ;
        END
    END IN
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 27.11  LAYER ME1  ;
        ANTENNADIFFAREA 21.33  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  16.22 1.90 16.50 2.50 ;
        RECT  16.22 0.64 16.50 1.24 ;
        RECT  16.22 0.64 16.38 2.50 ;
        RECT  0.74 1.52 16.38 1.68 ;
        RECT  15.18 1.90 15.46 2.50 ;
        RECT  15.18 0.64 15.46 1.24 ;
        RECT  15.24 0.64 15.40 2.50 ;
        RECT  14.14 1.90 14.42 2.50 ;
        RECT  14.14 0.64 14.42 1.24 ;
        RECT  14.20 0.64 14.36 2.50 ;
        RECT  13.10 1.90 13.38 2.50 ;
        RECT  13.10 0.64 13.38 1.24 ;
        RECT  13.16 0.64 13.32 2.50 ;
        RECT  12.06 1.90 12.34 2.50 ;
        RECT  12.06 0.64 12.34 1.24 ;
        RECT  12.12 0.64 12.28 2.50 ;
        RECT  11.02 1.90 11.30 2.50 ;
        RECT  11.02 0.64 11.30 1.24 ;
        RECT  11.08 0.64 11.24 2.50 ;
        RECT  9.98 1.90 10.26 2.50 ;
        RECT  9.98 0.64 10.26 1.24 ;
        RECT  10.04 0.64 10.20 2.50 ;
        RECT  8.94 1.90 9.22 2.50 ;
        RECT  8.94 0.64 9.22 1.24 ;
        RECT  9.00 0.64 9.16 2.50 ;
        RECT  7.90 1.90 8.18 2.50 ;
        RECT  7.90 0.64 8.18 1.24 ;
        RECT  7.96 0.64 8.12 2.50 ;
        RECT  6.86 1.90 7.14 2.50 ;
        RECT  6.86 0.64 7.14 1.24 ;
        RECT  6.92 0.64 7.08 2.50 ;
        RECT  5.82 1.90 6.10 2.50 ;
        RECT  5.82 0.64 6.10 1.24 ;
        RECT  5.88 0.64 6.04 2.50 ;
        RECT  4.78 1.90 5.06 2.50 ;
        RECT  4.78 0.64 5.06 1.24 ;
        RECT  4.84 0.64 5.00 2.50 ;
        RECT  3.74 1.90 4.02 2.50 ;
        RECT  3.74 0.64 4.02 1.24 ;
        RECT  3.80 0.64 3.96 2.50 ;
        RECT  2.70 1.90 2.98 2.50 ;
        RECT  2.70 0.64 2.98 1.24 ;
        RECT  2.76 0.64 2.92 2.50 ;
        RECT  1.66 1.90 1.94 2.50 ;
        RECT  1.66 0.64 1.94 1.24 ;
        RECT  1.72 0.64 1.88 2.50 ;
        RECT  0.74 1.46 1.14 1.74 ;
        RECT  0.62 1.90 0.90 2.50 ;
        RECT  0.74 0.64 0.90 2.50 ;
        RECT  0.62 0.64 0.90 1.24 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 17.20 3.48 ;
        RECT  16.74 2.88 17.02 3.48 ;
        RECT  16.74 1.90 17.02 2.50 ;
        RECT  16.80 1.90 16.96 3.48 ;
        RECT  15.70 1.90 15.98 2.50 ;
        RECT  15.76 1.90 15.92 3.48 ;
        RECT  14.66 1.90 14.94 2.50 ;
        RECT  14.72 1.90 14.88 3.48 ;
        RECT  13.62 1.90 13.90 2.50 ;
        RECT  13.68 1.90 13.84 3.48 ;
        RECT  12.58 1.90 12.86 2.50 ;
        RECT  12.64 1.90 12.80 3.48 ;
        RECT  11.54 1.90 11.82 2.50 ;
        RECT  11.60 1.90 11.76 3.48 ;
        RECT  10.50 1.90 10.78 2.50 ;
        RECT  10.56 1.90 10.72 3.48 ;
        RECT  9.46 1.90 9.74 2.50 ;
        RECT  9.52 1.90 9.68 3.48 ;
        RECT  8.42 1.90 8.70 2.50 ;
        RECT  8.48 1.90 8.64 3.48 ;
        RECT  7.38 1.90 7.66 2.50 ;
        RECT  7.44 1.90 7.60 3.48 ;
        RECT  6.34 1.90 6.62 2.50 ;
        RECT  6.40 1.90 6.56 3.48 ;
        RECT  5.30 1.90 5.58 2.50 ;
        RECT  5.36 1.90 5.52 3.48 ;
        RECT  4.26 1.90 4.54 2.50 ;
        RECT  4.32 1.90 4.48 3.48 ;
        RECT  3.22 1.90 3.50 2.50 ;
        RECT  3.28 1.90 3.44 3.48 ;
        RECT  2.18 1.90 2.46 2.50 ;
        RECT  2.24 1.90 2.40 3.48 ;
        RECT  1.14 1.90 1.42 2.50 ;
        RECT  1.20 1.90 1.36 3.48 ;
        RECT  0.10 1.90 0.38 2.50 ;
        RECT  0.16 1.90 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 17.20 0.28 ;
        RECT  16.74 0.64 17.02 1.24 ;
        RECT  16.74 -0.28 17.02 0.32 ;
        RECT  16.80 -0.28 16.96 1.24 ;
        RECT  15.70 0.64 15.98 1.24 ;
        RECT  15.76 -0.28 15.92 1.24 ;
        RECT  14.66 0.64 14.94 1.24 ;
        RECT  14.72 -0.28 14.88 1.24 ;
        RECT  13.62 0.64 13.90 1.24 ;
        RECT  13.68 -0.28 13.84 1.24 ;
        RECT  12.58 0.64 12.86 1.24 ;
        RECT  12.64 -0.28 12.80 1.24 ;
        RECT  11.54 0.64 11.82 1.24 ;
        RECT  11.60 -0.28 11.76 1.24 ;
        RECT  10.50 0.64 10.78 1.24 ;
        RECT  10.56 -0.28 10.72 1.24 ;
        RECT  9.46 0.64 9.74 1.24 ;
        RECT  9.52 -0.28 9.68 1.24 ;
        RECT  8.42 0.64 8.70 1.24 ;
        RECT  8.48 -0.28 8.64 1.24 ;
        RECT  7.38 0.64 7.66 1.24 ;
        RECT  7.44 -0.28 7.60 1.24 ;
        RECT  6.34 0.64 6.62 1.24 ;
        RECT  6.40 -0.28 6.56 1.24 ;
        RECT  5.30 0.64 5.58 1.24 ;
        RECT  5.36 -0.28 5.52 1.24 ;
        RECT  4.26 0.64 4.54 1.24 ;
        RECT  4.32 -0.28 4.48 1.24 ;
        RECT  3.22 0.64 3.50 1.24 ;
        RECT  3.28 -0.28 3.44 1.24 ;
        RECT  2.18 0.64 2.46 1.24 ;
        RECT  2.24 -0.28 2.40 1.24 ;
        RECT  1.14 0.64 1.42 1.24 ;
        RECT  1.20 -0.28 1.36 1.24 ;
        RECT  0.10 0.64 0.38 1.24 ;
        RECT  0.16 -0.28 0.32 1.24 ;
        END
    END GND!
END INVSP64V1_0

MACRO INVSP4V1_0
    CLASS CORE ;
    FOREIGN INVSP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 1.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 2.72  LAYER ME1  ;
        ANTENNADIFFAREA 1.94  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.82 1.46 1.14 1.74 ;
        RECT  0.70 1.90 0.98 2.50 ;
        RECT  0.82 0.64 0.98 2.50 ;
        RECT  0.70 0.64 0.98 1.24 ;
        END
    END OUT
    PIN IN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.29  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.46 0.64 1.74 ;
        END
    END IN
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 1.60 3.48 ;
        RECT  1.22 1.90 1.50 2.50 ;
        RECT  1.14 2.88 1.44 3.48 ;
        RECT  1.28 1.90 1.44 3.48 ;
        RECT  0.18 1.90 0.46 2.50 ;
        RECT  0.24 1.90 0.40 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 1.60 0.28 ;
        RECT  1.22 0.64 1.50 1.24 ;
        RECT  1.28 -0.28 1.44 1.24 ;
        RECT  1.14 -0.28 1.44 0.32 ;
        RECT  0.18 0.64 0.46 1.24 ;
        RECT  0.24 -0.28 0.40 1.24 ;
        END
    END GND!
END INVSP4V1_0

MACRO INVSP48V1_0
    CLASS CORE ;
    FOREIGN INVSP48V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 13.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 3.46  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.46 0.56 1.74 ;
        END
    END IN
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 20.79  LAYER ME1  ;
        ANTENNADIFFAREA 16.21  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.06 1.90 12.34 2.50 ;
        RECT  12.06 0.64 12.34 1.24 ;
        RECT  12.06 0.64 12.22 2.50 ;
        RECT  0.74 1.52 12.22 1.68 ;
        RECT  11.02 1.90 11.30 2.50 ;
        RECT  11.02 0.64 11.30 1.24 ;
        RECT  11.08 0.64 11.24 2.50 ;
        RECT  9.98 1.90 10.26 2.50 ;
        RECT  9.98 0.64 10.26 1.24 ;
        RECT  10.04 0.64 10.20 2.50 ;
        RECT  8.94 1.90 9.22 2.50 ;
        RECT  8.94 0.64 9.22 1.24 ;
        RECT  9.00 0.64 9.16 2.50 ;
        RECT  7.90 1.90 8.18 2.50 ;
        RECT  7.90 0.64 8.18 1.24 ;
        RECT  7.96 0.64 8.12 2.50 ;
        RECT  6.86 1.90 7.14 2.50 ;
        RECT  6.86 0.64 7.14 1.24 ;
        RECT  6.92 0.64 7.08 2.50 ;
        RECT  5.82 1.90 6.10 2.50 ;
        RECT  5.82 0.64 6.10 1.24 ;
        RECT  5.88 0.64 6.04 2.50 ;
        RECT  4.78 1.90 5.06 2.50 ;
        RECT  4.78 0.64 5.06 1.24 ;
        RECT  4.84 0.64 5.00 2.50 ;
        RECT  3.74 1.90 4.02 2.50 ;
        RECT  3.74 0.64 4.02 1.24 ;
        RECT  3.80 0.64 3.96 2.50 ;
        RECT  2.70 1.90 2.98 2.50 ;
        RECT  2.70 0.64 2.98 1.24 ;
        RECT  2.76 0.64 2.92 2.50 ;
        RECT  1.66 1.90 1.94 2.50 ;
        RECT  1.66 0.64 1.94 1.24 ;
        RECT  1.72 0.64 1.88 2.50 ;
        RECT  0.74 1.46 1.14 1.74 ;
        RECT  0.62 1.90 0.90 2.50 ;
        RECT  0.74 0.64 0.90 2.50 ;
        RECT  0.62 0.64 0.90 1.24 ;
        END
    END OUT
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 13.20 0.28 ;
        RECT  12.64 -0.28 13.02 0.32 ;
        RECT  12.58 0.64 12.86 1.24 ;
        RECT  12.64 -0.28 12.80 1.24 ;
        RECT  11.54 0.64 11.82 1.24 ;
        RECT  11.60 -0.28 11.76 1.24 ;
        RECT  10.50 0.64 10.78 1.24 ;
        RECT  10.56 -0.28 10.72 1.24 ;
        RECT  9.46 0.64 9.74 1.24 ;
        RECT  9.52 -0.28 9.68 1.24 ;
        RECT  8.42 0.64 8.70 1.24 ;
        RECT  8.48 -0.28 8.64 1.24 ;
        RECT  7.38 0.64 7.66 1.24 ;
        RECT  7.44 -0.28 7.60 1.24 ;
        RECT  6.34 0.64 6.62 1.24 ;
        RECT  6.40 -0.28 6.56 1.24 ;
        RECT  5.30 0.64 5.58 1.24 ;
        RECT  5.36 -0.28 5.52 1.24 ;
        RECT  4.26 0.64 4.54 1.24 ;
        RECT  4.32 -0.28 4.48 1.24 ;
        RECT  3.22 0.64 3.50 1.24 ;
        RECT  3.28 -0.28 3.44 1.24 ;
        RECT  2.18 0.64 2.46 1.24 ;
        RECT  2.24 -0.28 2.40 1.24 ;
        RECT  1.14 0.64 1.42 1.24 ;
        RECT  1.20 -0.28 1.36 1.24 ;
        RECT  0.10 0.64 0.38 1.24 ;
        RECT  0.16 -0.28 0.32 1.24 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 13.20 3.48 ;
        RECT  12.64 2.88 13.02 3.48 ;
        RECT  12.58 1.90 12.86 2.50 ;
        RECT  12.64 1.90 12.80 3.48 ;
        RECT  11.54 1.90 11.82 2.50 ;
        RECT  11.60 1.90 11.76 3.48 ;
        RECT  10.50 1.90 10.78 2.50 ;
        RECT  10.56 1.90 10.72 3.48 ;
        RECT  9.46 1.90 9.74 2.50 ;
        RECT  9.52 1.90 9.68 3.48 ;
        RECT  8.42 1.90 8.70 2.50 ;
        RECT  8.48 1.90 8.64 3.48 ;
        RECT  7.38 1.90 7.66 2.50 ;
        RECT  7.44 1.90 7.60 3.48 ;
        RECT  6.34 1.90 6.62 2.50 ;
        RECT  6.40 1.90 6.56 3.48 ;
        RECT  5.30 1.90 5.58 2.50 ;
        RECT  5.36 1.90 5.52 3.48 ;
        RECT  4.26 1.90 4.54 2.50 ;
        RECT  4.32 1.90 4.48 3.48 ;
        RECT  3.22 1.90 3.50 2.50 ;
        RECT  3.28 1.90 3.44 3.48 ;
        RECT  2.18 1.90 2.46 2.50 ;
        RECT  2.24 1.90 2.40 3.48 ;
        RECT  1.14 1.90 1.42 2.50 ;
        RECT  1.20 1.90 1.36 3.48 ;
        RECT  0.10 1.90 0.38 2.50 ;
        RECT  0.16 1.90 0.32 3.48 ;
        END
    END VDD!
END INVSP48V1_0

MACRO INVSP32V1_0
    CLASS CORE ;
    FOREIGN INVSP32V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.30  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.46 0.56 1.74 ;
        END
    END IN
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 14.01  LAYER ME1  ;
        ANTENNADIFFAREA 10.97  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.90 1.90 8.18 2.50 ;
        RECT  7.90 0.64 8.18 1.24 ;
        RECT  7.90 0.64 8.06 2.50 ;
        RECT  0.74 1.52 8.06 1.68 ;
        RECT  6.86 1.90 7.14 2.50 ;
        RECT  6.86 0.64 7.14 1.24 ;
        RECT  6.92 0.64 7.08 2.50 ;
        RECT  5.82 1.90 6.10 2.50 ;
        RECT  5.82 0.64 6.10 1.24 ;
        RECT  5.88 0.64 6.04 2.50 ;
        RECT  4.78 1.90 5.06 2.50 ;
        RECT  4.78 0.64 5.06 1.24 ;
        RECT  4.84 0.64 5.00 2.50 ;
        RECT  3.74 1.90 4.02 2.50 ;
        RECT  3.74 0.64 4.02 1.24 ;
        RECT  3.80 0.64 3.96 2.50 ;
        RECT  2.70 1.90 2.98 2.50 ;
        RECT  2.70 0.64 2.98 1.24 ;
        RECT  2.76 0.64 2.92 2.50 ;
        RECT  1.66 1.90 1.94 2.50 ;
        RECT  1.66 0.64 1.94 1.24 ;
        RECT  1.72 0.64 1.88 2.50 ;
        RECT  0.74 1.46 1.14 1.74 ;
        RECT  0.62 1.90 0.90 2.50 ;
        RECT  0.74 0.64 0.90 2.50 ;
        RECT  0.62 0.64 0.90 1.24 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 8.80 3.48 ;
        RECT  8.42 1.90 8.70 2.50 ;
        RECT  8.34 2.88 8.64 3.48 ;
        RECT  8.48 1.90 8.64 3.48 ;
        RECT  7.38 1.90 7.66 2.50 ;
        RECT  7.44 1.90 7.60 3.48 ;
        RECT  6.34 1.90 6.62 2.50 ;
        RECT  6.40 1.90 6.56 3.48 ;
        RECT  5.30 1.90 5.58 2.50 ;
        RECT  5.36 1.90 5.52 3.48 ;
        RECT  4.26 1.90 4.54 2.50 ;
        RECT  4.32 1.90 4.48 3.48 ;
        RECT  3.22 1.90 3.50 2.50 ;
        RECT  3.28 1.90 3.44 3.48 ;
        RECT  2.18 1.90 2.46 2.50 ;
        RECT  2.24 1.90 2.40 3.48 ;
        RECT  1.14 1.90 1.42 2.50 ;
        RECT  1.20 1.90 1.36 3.48 ;
        RECT  0.10 1.90 0.38 2.50 ;
        RECT  0.16 1.90 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 8.80 0.28 ;
        RECT  8.42 0.64 8.70 1.24 ;
        RECT  8.48 -0.28 8.64 1.24 ;
        RECT  8.34 -0.28 8.64 0.32 ;
        RECT  7.38 0.64 7.66 1.24 ;
        RECT  7.44 -0.28 7.60 1.24 ;
        RECT  6.34 0.64 6.62 1.24 ;
        RECT  6.40 -0.28 6.56 1.24 ;
        RECT  5.30 0.64 5.58 1.24 ;
        RECT  5.36 -0.28 5.52 1.24 ;
        RECT  4.26 0.64 4.54 1.24 ;
        RECT  4.32 -0.28 4.48 1.24 ;
        RECT  3.22 0.64 3.50 1.24 ;
        RECT  3.28 -0.28 3.44 1.24 ;
        RECT  2.18 0.64 2.46 1.24 ;
        RECT  2.24 -0.28 2.40 1.24 ;
        RECT  1.14 0.64 1.42 1.24 ;
        RECT  1.20 -0.28 1.36 1.24 ;
        RECT  0.10 0.64 0.38 1.24 ;
        RECT  0.16 -0.28 0.32 1.24 ;
        END
    END GND!
END INVSP32V1_0

MACRO INVSP2V1_0
    CLASS CORE ;
    FOREIGN INVSP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 1.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.14  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.44 1.46 0.86 1.74 ;
        END
    END IN
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 1.82  LAYER ME1  ;
        ANTENNADIFFAREA 1.33  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.90 0.38 2.50 ;
        RECT  0.10 0.64 0.38 1.24 ;
        RECT  0.12 0.64 0.28 2.50 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 1.20 3.48 ;
        RECT  0.68 2.88 1.02 3.48 ;
        RECT  0.62 1.90 0.90 2.50 ;
        RECT  0.68 1.90 0.84 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 1.20 0.28 ;
        RECT  0.68 -0.28 1.02 0.32 ;
        RECT  0.62 0.64 0.90 1.24 ;
        RECT  0.68 -0.28 0.84 1.24 ;
        END
    END GND!
END INVSP2V1_0

MACRO INVSP24V1_0
    CLASS CORE ;
    FOREIGN INVSP24V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.73  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.46 0.56 1.74 ;
        END
    END IN
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 10.85  LAYER ME1  ;
        ANTENNADIFFAREA 8.41  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.82 1.90 6.10 2.50 ;
        RECT  5.82 0.64 6.10 1.24 ;
        RECT  5.82 0.64 5.98 2.50 ;
        RECT  0.74 1.52 5.98 1.68 ;
        RECT  4.78 1.90 5.06 2.50 ;
        RECT  4.78 0.64 5.06 1.24 ;
        RECT  4.84 0.64 5.00 2.50 ;
        RECT  3.74 1.90 4.02 2.50 ;
        RECT  3.74 0.64 4.02 1.24 ;
        RECT  3.80 0.64 3.96 2.50 ;
        RECT  2.70 1.90 2.98 2.50 ;
        RECT  2.70 0.64 2.98 1.24 ;
        RECT  2.76 0.64 2.92 2.50 ;
        RECT  1.66 1.90 1.94 2.50 ;
        RECT  1.66 0.64 1.94 1.24 ;
        RECT  1.72 0.64 1.88 2.50 ;
        RECT  0.74 1.46 1.14 1.74 ;
        RECT  0.62 1.90 0.90 2.50 ;
        RECT  0.74 0.64 0.90 2.50 ;
        RECT  0.62 0.64 0.90 1.24 ;
        END
    END OUT
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 6.80 0.28 ;
        RECT  6.34 0.64 6.62 1.24 ;
        RECT  6.34 -0.28 6.62 0.32 ;
        RECT  6.40 -0.28 6.56 1.24 ;
        RECT  5.30 0.64 5.58 1.24 ;
        RECT  5.36 -0.28 5.52 1.24 ;
        RECT  4.26 0.64 4.54 1.24 ;
        RECT  4.32 -0.28 4.48 1.24 ;
        RECT  3.22 0.64 3.50 1.24 ;
        RECT  3.28 -0.28 3.44 1.24 ;
        RECT  2.18 0.64 2.46 1.24 ;
        RECT  2.24 -0.28 2.40 1.24 ;
        RECT  1.14 0.64 1.42 1.24 ;
        RECT  1.20 -0.28 1.36 1.24 ;
        RECT  0.10 0.64 0.38 1.24 ;
        RECT  0.16 -0.28 0.32 1.24 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 6.80 3.48 ;
        RECT  6.34 2.88 6.62 3.48 ;
        RECT  6.34 1.90 6.62 2.50 ;
        RECT  6.40 1.90 6.56 3.48 ;
        RECT  5.30 1.90 5.58 2.50 ;
        RECT  5.36 1.90 5.52 3.48 ;
        RECT  4.26 1.90 4.54 2.50 ;
        RECT  4.32 1.90 4.48 3.48 ;
        RECT  3.22 1.90 3.50 2.50 ;
        RECT  3.28 1.90 3.44 3.48 ;
        RECT  2.18 1.90 2.46 2.50 ;
        RECT  2.24 1.90 2.40 3.48 ;
        RECT  1.14 1.90 1.42 2.50 ;
        RECT  1.20 1.90 1.36 3.48 ;
        RECT  0.10 1.90 0.38 2.50 ;
        RECT  0.16 1.90 0.32 3.48 ;
        END
    END VDD!
END INVSP24V1_0

MACRO INVSP1V1_0
    CLASS CORE ;
    FOREIGN INVSP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 1.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.44 1.46 0.86 1.74 ;
        END
    END IN
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 1.74  LAYER ME1  ;
        ANTENNADIFFAREA 0.90  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.12 1.90 0.40 2.18 ;
        RECT  0.12 0.96 0.40 1.24 ;
        RECT  0.12 0.96 0.28 2.18 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 1.20 3.48 ;
        RECT  0.70 2.88 1.02 3.48 ;
        RECT  0.64 1.90 0.92 2.18 ;
        RECT  0.70 1.90 0.86 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 1.20 0.28 ;
        RECT  0.70 -0.28 1.02 0.32 ;
        RECT  0.64 0.96 0.92 1.24 ;
        RECT  0.70 -0.28 0.86 1.24 ;
        END
    END GND!
END INVSP1V1_0

MACRO INVSP16V1_0
    CLASS CORE ;
    FOREIGN INVSP16V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.46 0.56 1.74 ;
        END
    END IN
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 7.69  LAYER ME1  ;
        ANTENNADIFFAREA 5.85  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.74 1.90 4.02 2.50 ;
        RECT  3.74 0.64 4.02 1.24 ;
        RECT  3.74 0.64 3.90 2.50 ;
        RECT  0.74 1.52 3.90 1.68 ;
        RECT  2.70 1.90 2.98 2.50 ;
        RECT  2.70 0.64 2.98 1.24 ;
        RECT  2.76 0.64 2.92 2.50 ;
        RECT  1.66 1.90 1.94 2.50 ;
        RECT  1.66 0.64 1.94 1.24 ;
        RECT  1.72 0.64 1.88 2.50 ;
        RECT  0.74 1.46 1.14 1.74 ;
        RECT  0.62 1.90 0.90 2.50 ;
        RECT  0.74 0.64 0.90 2.50 ;
        RECT  0.62 0.64 0.90 1.24 ;
        END
    END OUT
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.80 0.28 ;
        RECT  4.32 -0.28 4.62 0.32 ;
        RECT  4.26 0.64 4.54 1.24 ;
        RECT  4.32 -0.28 4.48 1.24 ;
        RECT  3.22 0.64 3.50 1.24 ;
        RECT  3.28 -0.28 3.44 1.24 ;
        RECT  2.18 0.64 2.46 1.24 ;
        RECT  2.24 -0.28 2.40 1.24 ;
        RECT  1.14 0.64 1.42 1.24 ;
        RECT  1.20 -0.28 1.36 1.24 ;
        RECT  0.10 0.64 0.38 1.24 ;
        RECT  0.16 -0.28 0.32 1.24 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.80 3.48 ;
        RECT  4.32 2.88 4.62 3.48 ;
        RECT  4.26 1.90 4.54 2.50 ;
        RECT  4.32 1.90 4.48 3.48 ;
        RECT  3.22 1.90 3.50 2.50 ;
        RECT  3.28 1.90 3.44 3.48 ;
        RECT  2.18 1.90 2.46 2.50 ;
        RECT  2.24 1.90 2.40 3.48 ;
        RECT  1.14 1.90 1.42 2.50 ;
        RECT  1.20 1.90 1.36 3.48 ;
        RECT  0.10 1.90 0.38 2.50 ;
        RECT  0.16 1.90 0.32 3.48 ;
        END
    END VDD!
END INVSP16V1_0

MACRO INVSP12V1_0
    CLASS CORE ;
    FOREIGN INVSP12V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.86  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.46 0.56 1.74 ;
        END
    END IN
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 5.89  LAYER ME1  ;
        ANTENNADIFFAREA 4.50  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.70 1.90 2.98 2.50 ;
        RECT  2.70 0.64 2.98 1.24 ;
        RECT  2.70 0.64 2.86 2.50 ;
        RECT  0.74 1.52 2.86 1.68 ;
        RECT  1.66 1.90 1.94 2.50 ;
        RECT  1.66 0.64 1.94 1.24 ;
        RECT  1.72 0.64 1.88 2.50 ;
        RECT  0.74 1.46 1.14 1.74 ;
        RECT  0.62 1.90 0.90 2.50 ;
        RECT  0.74 0.64 0.90 2.50 ;
        RECT  0.62 0.64 0.90 1.24 ;
        END
    END OUT
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 3.60 0.28 ;
        RECT  3.22 0.64 3.50 1.24 ;
        RECT  3.28 -0.28 3.44 1.24 ;
        RECT  3.14 -0.28 3.44 0.32 ;
        RECT  2.18 0.64 2.46 1.24 ;
        RECT  2.24 -0.28 2.40 1.24 ;
        RECT  1.14 0.64 1.42 1.24 ;
        RECT  1.20 -0.28 1.36 1.24 ;
        RECT  0.10 0.64 0.38 1.24 ;
        RECT  0.16 -0.28 0.32 1.24 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 3.60 3.48 ;
        RECT  3.22 1.90 3.50 2.50 ;
        RECT  3.14 2.88 3.44 3.48 ;
        RECT  3.28 1.90 3.44 3.48 ;
        RECT  2.18 1.90 2.46 2.50 ;
        RECT  2.24 1.90 2.40 3.48 ;
        RECT  1.14 1.90 1.42 2.50 ;
        RECT  1.20 1.90 1.36 3.48 ;
        RECT  0.10 1.90 0.38 2.50 ;
        RECT  0.16 1.90 0.32 3.48 ;
        END
    END VDD!
END INVSP12V1_0

MACRO INVCKSP8V1_0
    CLASS CORE ;
    FOREIGN INVCKSP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.75  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.79 1.06 3.21 1.34 ;
        END
    END IN
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 6.17  LAYER ME1  ;
        ANTENNADIFFAREA 4.26  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.70 1.84 2.98 2.62 ;
        RECT  2.70 1.52 2.86 2.62 ;
        RECT  0.74 1.52 2.86 1.68 ;
        RECT  1.66 1.84 1.94 2.62 ;
        RECT  1.66 0.84 1.94 1.24 ;
        RECT  1.72 0.84 1.88 2.62 ;
        RECT  0.62 1.84 0.90 2.62 ;
        RECT  0.74 0.84 0.90 2.62 ;
        RECT  0.62 0.84 0.90 1.24 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.00 3.48 ;
        RECT  3.54 2.88 3.82 3.48 ;
        RECT  3.22 1.84 3.50 2.62 ;
        RECT  3.22 1.84 3.38 3.48 ;
        RECT  2.18 1.84 2.46 2.62 ;
        RECT  2.24 1.84 2.40 3.48 ;
        RECT  1.14 1.84 1.42 2.62 ;
        RECT  1.20 1.84 1.36 3.48 ;
        RECT  0.10 1.84 0.38 2.62 ;
        RECT  0.16 1.84 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.00 0.28 ;
        RECT  3.54 -0.28 3.82 0.32 ;
        RECT  2.18 0.84 2.46 1.24 ;
        RECT  2.24 -0.28 2.40 1.24 ;
        RECT  1.14 0.84 1.42 1.24 ;
        RECT  1.20 -0.28 1.36 1.24 ;
        RECT  0.10 0.84 0.38 1.24 ;
        RECT  0.16 -0.28 0.32 1.24 ;
        END
    END GND!
END INVCKSP8V1_0

MACRO INVCKSP4V1_0
    CLASS CORE ;
    FOREIGN INVCKSP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 2.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 3.65  LAYER ME1  ;
        ANTENNADIFFAREA 2.54  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.66 1.86 1.94 2.66 ;
        RECT  1.66 1.48 1.82 2.66 ;
        RECT  0.74 1.48 1.82 1.64 ;
        RECT  0.62 1.86 0.90 2.66 ;
        RECT  0.74 0.82 0.90 2.66 ;
        RECT  0.62 0.82 0.90 1.24 ;
        END
    END OUT
    PIN IN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.39  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.06 1.36 2.32 1.74 ;
        RECT  2.02 1.44 2.32 1.72 ;
        END
    END IN
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 2.40 3.48 ;
        RECT  1.94 2.88 2.22 3.48 ;
        RECT  1.14 1.86 1.42 2.66 ;
        RECT  1.20 1.86 1.36 3.48 ;
        RECT  0.10 1.86 0.38 2.66 ;
        RECT  0.16 1.86 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 2.40 0.28 ;
        RECT  1.94 -0.28 2.22 0.32 ;
        RECT  1.14 0.82 1.42 1.24 ;
        RECT  1.20 -0.28 1.36 1.24 ;
        RECT  0.10 0.82 0.38 1.24 ;
        RECT  0.16 -0.28 0.32 1.24 ;
        END
    END GND!
END INVCKSP4V1_0

MACRO INVCKSP32V1_0
    CLASS CORE ;
    FOREIGN INVCKSP32V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 13.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 3.08  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.39 1.06 0.81 1.34 ;
        END
    END IN
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 19.97  LAYER ME1  ;
        ANTENNADIFFAREA 14.97  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.06 1.84 12.34 2.64 ;
        RECT  12.06 1.52 12.22 2.64 ;
        RECT  0.74 1.52 12.22 1.68 ;
        RECT  11.02 1.84 11.30 2.64 ;
        RECT  11.08 1.52 11.24 2.64 ;
        RECT  9.98 1.84 10.26 2.64 ;
        RECT  10.04 1.52 10.20 2.64 ;
        RECT  9.46 0.78 9.74 1.24 ;
        RECT  9.52 0.78 9.68 1.68 ;
        RECT  8.94 1.84 9.22 2.64 ;
        RECT  9.00 1.52 9.16 2.64 ;
        RECT  8.42 0.78 8.70 1.24 ;
        RECT  8.48 0.78 8.64 1.68 ;
        RECT  7.90 1.84 8.18 2.64 ;
        RECT  7.96 1.52 8.12 2.64 ;
        RECT  7.38 0.78 7.66 1.24 ;
        RECT  7.44 0.78 7.60 1.68 ;
        RECT  6.86 1.84 7.14 2.64 ;
        RECT  6.92 1.52 7.08 2.64 ;
        RECT  6.34 0.78 6.62 1.24 ;
        RECT  6.40 0.78 6.56 1.68 ;
        RECT  5.82 1.84 6.10 2.64 ;
        RECT  5.88 1.52 6.04 2.64 ;
        RECT  5.30 0.78 5.58 1.24 ;
        RECT  5.36 0.78 5.52 1.68 ;
        RECT  4.78 1.84 5.06 2.64 ;
        RECT  4.84 1.52 5.00 2.64 ;
        RECT  4.26 0.78 4.54 1.24 ;
        RECT  4.32 0.78 4.48 1.68 ;
        RECT  3.74 1.84 4.02 2.64 ;
        RECT  3.80 1.52 3.96 2.64 ;
        RECT  3.22 0.78 3.50 1.24 ;
        RECT  3.28 0.78 3.44 1.68 ;
        RECT  2.70 1.84 2.98 2.64 ;
        RECT  2.76 1.52 2.92 2.64 ;
        RECT  1.66 1.84 1.94 2.64 ;
        RECT  1.72 1.52 1.88 2.64 ;
        RECT  0.62 1.84 0.90 2.64 ;
        RECT  0.74 1.52 0.90 2.64 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 13.20 3.48 ;
        RECT  12.64 2.88 13.02 3.48 ;
        RECT  12.58 1.84 12.86 2.64 ;
        RECT  12.64 1.84 12.80 3.48 ;
        RECT  11.54 1.84 11.82 2.64 ;
        RECT  11.60 1.84 11.76 3.48 ;
        RECT  10.50 1.84 10.78 2.64 ;
        RECT  10.56 1.84 10.72 3.48 ;
        RECT  9.46 1.84 9.74 2.64 ;
        RECT  9.52 1.84 9.68 3.48 ;
        RECT  8.42 1.84 8.70 2.64 ;
        RECT  8.48 1.84 8.64 3.48 ;
        RECT  7.38 1.84 7.66 2.64 ;
        RECT  7.44 1.84 7.60 3.48 ;
        RECT  6.34 1.84 6.62 2.64 ;
        RECT  6.40 1.84 6.56 3.48 ;
        RECT  5.30 1.84 5.58 2.64 ;
        RECT  5.36 1.84 5.52 3.48 ;
        RECT  4.26 1.84 4.54 2.64 ;
        RECT  4.32 1.84 4.48 3.48 ;
        RECT  3.22 1.84 3.50 2.64 ;
        RECT  3.28 1.84 3.44 3.48 ;
        RECT  2.18 1.84 2.46 2.64 ;
        RECT  2.24 1.84 2.40 3.48 ;
        RECT  1.14 1.84 1.42 2.64 ;
        RECT  1.20 1.84 1.36 3.48 ;
        RECT  0.10 1.84 0.38 2.64 ;
        RECT  0.16 1.84 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 13.20 0.28 ;
        RECT  12.74 -0.28 13.02 0.32 ;
        RECT  9.98 0.78 10.26 1.24 ;
        RECT  10.04 -0.28 10.20 1.24 ;
        RECT  8.94 0.78 9.22 1.24 ;
        RECT  9.00 -0.28 9.16 1.24 ;
        RECT  7.90 0.78 8.18 1.24 ;
        RECT  7.96 -0.28 8.12 1.24 ;
        RECT  6.86 0.78 7.14 1.24 ;
        RECT  6.92 -0.28 7.08 1.24 ;
        RECT  5.82 0.78 6.10 1.24 ;
        RECT  5.88 -0.28 6.04 1.24 ;
        RECT  4.78 0.78 5.06 1.24 ;
        RECT  4.84 -0.28 5.00 1.24 ;
        RECT  3.74 0.78 4.02 1.24 ;
        RECT  3.80 -0.28 3.96 1.24 ;
        RECT  2.70 0.78 2.98 1.24 ;
        RECT  2.76 -0.28 2.92 1.24 ;
        END
    END GND!
END INVCKSP32V1_0

MACRO INVCKSP2V1_0
    CLASS CORE ;
    FOREIGN INVCKSP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 1.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.16  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.46 0.49 1.74 ;
        END
    END IN
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 2.45  LAYER ME1  ;
        ANTENNADIFFAREA 1.43  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.78 1.46 1.14 1.74 ;
        RECT  0.66 1.90 0.94 2.42 ;
        RECT  0.78 0.92 0.94 2.42 ;
        RECT  0.66 0.92 0.94 1.24 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 1.60 3.48 ;
        RECT  1.18 1.90 1.46 2.42 ;
        RECT  1.14 2.88 1.42 3.48 ;
        RECT  1.24 1.90 1.40 3.48 ;
        RECT  0.14 1.90 0.42 2.42 ;
        RECT  0.20 1.90 0.36 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 1.60 0.28 ;
        RECT  1.14 -0.28 1.42 0.32 ;
        RECT  0.14 0.92 0.42 1.24 ;
        RECT  0.20 -0.28 0.36 1.24 ;
        END
    END GND!
END INVCKSP2V1_0

MACRO INVCKSP1V1_0
    CLASS CORE ;
    FOREIGN INVCKSP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 1.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 1.78  LAYER ME1  ;
        ANTENNADIFFAREA 1.14  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.12 1.90 0.42 2.54 ;
        RECT  0.10 0.96 0.38 1.24 ;
        RECT  0.12 0.96 0.28 2.54 ;
        END
    END OUT
    PIN IN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.10  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.44 1.46 0.86 1.74 ;
        END
    END IN
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 1.20 3.48 ;
        RECT  0.72 2.88 1.02 3.48 ;
        RECT  0.66 1.90 0.94 2.54 ;
        RECT  0.72 1.90 0.88 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 1.20 0.28 ;
        RECT  0.72 -0.28 1.02 0.32 ;
        RECT  0.70 0.96 0.98 1.24 ;
        RECT  0.72 -0.28 0.88 1.24 ;
        END
    END GND!
END INVCKSP1V1_0

MACRO INVCKSP16V1_0
    CLASS CORE ;
    FOREIGN INVCKSP16V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.54  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.39 1.06 0.81 1.34 ;
        END
    END IN
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 10.80  LAYER ME1  ;
        ANTENNADIFFAREA 7.92  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.82 1.84 6.10 2.64 ;
        RECT  5.88 1.52 6.04 2.64 ;
        RECT  0.74 1.52 6.04 1.68 ;
        RECT  4.78 1.84 5.06 2.64 ;
        RECT  4.78 0.78 5.06 1.24 ;
        RECT  4.84 0.78 5.00 2.64 ;
        RECT  3.74 1.84 4.02 2.64 ;
        RECT  3.74 0.78 4.02 1.24 ;
        RECT  3.80 0.78 3.96 2.64 ;
        RECT  2.70 1.84 2.98 2.64 ;
        RECT  2.70 0.78 2.98 1.24 ;
        RECT  2.76 0.78 2.92 2.64 ;
        RECT  1.66 1.84 1.94 2.64 ;
        RECT  1.66 0.78 1.94 1.24 ;
        RECT  1.72 0.78 1.88 2.64 ;
        RECT  0.62 1.84 0.90 2.64 ;
        RECT  0.74 1.52 0.90 2.64 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 7.20 3.48 ;
        RECT  6.74 2.88 7.02 3.48 ;
        RECT  6.34 1.84 6.62 2.64 ;
        RECT  6.40 1.84 6.56 3.48 ;
        RECT  5.30 1.84 5.58 2.64 ;
        RECT  5.36 1.84 5.52 3.48 ;
        RECT  4.26 1.84 4.54 2.64 ;
        RECT  4.32 1.84 4.48 3.48 ;
        RECT  3.22 1.84 3.50 2.64 ;
        RECT  3.28 1.84 3.44 3.48 ;
        RECT  2.18 1.84 2.46 2.64 ;
        RECT  2.24 1.84 2.40 3.48 ;
        RECT  1.14 1.84 1.42 2.64 ;
        RECT  1.20 1.84 1.36 3.48 ;
        RECT  0.10 1.84 0.38 2.64 ;
        RECT  0.16 1.84 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 7.20 0.28 ;
        RECT  6.74 -0.28 7.02 0.32 ;
        RECT  4.26 0.78 4.54 1.24 ;
        RECT  4.32 -0.28 4.48 1.24 ;
        RECT  3.22 0.78 3.50 1.24 ;
        RECT  3.28 -0.28 3.44 1.24 ;
        RECT  2.18 0.78 2.46 1.24 ;
        RECT  2.24 -0.28 2.40 1.24 ;
        RECT  1.14 0.78 1.42 1.24 ;
        RECT  1.20 -0.28 1.36 1.24 ;
        END
    END GND!
END INVCKSP16V1_0

MACRO HASP8V1_0
    CLASS CORE ;
    FOREIGN HASP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN C
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 19.31  LAYER ME1  ;
        ANTENNADIFFAREA 10.09  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.29  LAYER ME1  ;
        ANTENNAMAXAREACAR 15.01  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.66 1.84 1.94 2.44 ;
        RECT  1.66 0.64 1.94 1.24 ;
        RECT  1.66 0.64 1.82 2.44 ;
        RECT  0.52 1.52 1.82 1.68 ;
        RECT  0.62 1.84 0.90 2.44 ;
        RECT  0.62 0.64 0.90 1.24 ;
        RECT  0.62 0.64 0.78 2.44 ;
        END
    END C
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 19.31  LAYER ME1  ;
        ANTENNADIFFAREA 10.09  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.29  LAYER ME1  ;
        ANTENNAMAXAREACAR 15.01  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.69 1.86 8.97 2.46 ;
        RECT  8.69 0.64 8.97 1.24 ;
        RECT  8.69 0.64 8.85 2.46 ;
        RECT  7.81 1.52 8.85 1.68 ;
        RECT  7.65 1.86 7.97 2.46 ;
        RECT  7.81 0.64 7.97 2.46 ;
        RECT  7.65 0.64 7.97 1.24 ;
        END
    END OUT
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.81 1.40 7.17 1.70 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.06 1.52 4.34 1.94 ;
        END
    END A
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 9.60 0.28 ;
        RECT  9.21 0.64 9.49 1.24 ;
        RECT  9.27 -0.28 9.43 1.24 ;
        RECT  9.14 -0.28 9.43 0.32 ;
        RECT  8.17 0.64 8.45 1.24 ;
        RECT  8.23 -0.28 8.39 1.24 ;
        RECT  7.13 0.64 7.41 1.24 ;
        RECT  7.19 -0.28 7.35 1.24 ;
        RECT  4.11 0.76 4.39 1.04 ;
        RECT  4.17 -0.28 4.33 1.04 ;
        RECT  2.18 0.64 2.46 1.24 ;
        RECT  2.24 -0.28 2.40 1.24 ;
        RECT  1.14 0.64 1.42 1.24 ;
        RECT  1.20 -0.28 1.36 1.24 ;
        RECT  0.10 0.64 0.38 1.24 ;
        RECT  0.16 -0.28 0.32 1.24 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 9.60 3.48 ;
        RECT  9.21 1.86 9.49 2.46 ;
        RECT  9.14 2.88 9.43 3.48 ;
        RECT  9.27 1.86 9.43 3.48 ;
        RECT  8.17 1.86 8.45 2.46 ;
        RECT  8.23 1.86 8.39 3.48 ;
        RECT  6.99 2.62 7.27 3.48 ;
        RECT  4.39 2.16 4.67 2.44 ;
        RECT  4.45 2.16 4.61 3.48 ;
        RECT  3.26 1.84 3.54 2.12 ;
        RECT  3.32 1.84 3.48 3.48 ;
        RECT  2.18 1.84 2.46 2.44 ;
        RECT  2.24 1.84 2.40 3.48 ;
        RECT  1.14 1.84 1.42 2.44 ;
        RECT  1.20 1.84 1.36 3.48 ;
        RECT  0.10 1.84 0.38 2.44 ;
        RECT  0.16 1.84 0.32 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  3.06 0.96 3.34 1.24 ;
        RECT  2.82 1.08 3.34 1.24 ;
        RECT  2.00 1.46 2.98 1.62 ;
        RECT  2.00 1.40 2.28 1.68 ;
        RECT  2.82 1.08 2.98 2.12 ;
        RECT  2.74 1.84 3.02 2.12 ;
        RECT  4.87 0.76 5.17 1.04 ;
        RECT  5.01 0.76 5.17 2.44 ;
        RECT  4.91 2.16 5.19 2.44 ;
        RECT  4.55 0.44 6.07 0.60 ;
        RECT  3.59 0.76 3.87 1.04 ;
        RECT  5.91 0.76 6.19 1.04 ;
        RECT  4.55 0.44 4.71 1.36 ;
        RECT  3.71 1.20 4.85 1.36 ;
        RECT  4.57 1.20 4.85 1.48 ;
        RECT  3.71 0.76 3.87 2.44 ;
        RECT  5.91 0.44 6.07 2.44 ;
        RECT  3.71 2.16 4.15 2.44 ;
        RECT  5.91 2.16 6.23 2.44 ;
        RECT  6.49 0.96 6.85 1.24 ;
        RECT  6.37 1.40 6.65 1.68 ;
        RECT  6.49 0.96 6.65 2.14 ;
        RECT  6.49 1.86 6.85 2.14 ;
        RECT  5.39 0.76 5.67 1.04 ;
        RECT  7.33 1.40 7.65 1.68 ;
        RECT  5.49 0.76 5.65 2.44 ;
        RECT  5.43 2.16 5.71 2.44 ;
        RECT  7.33 1.40 7.49 2.46 ;
        RECT  6.39 2.30 7.49 2.46 ;
        RECT  5.55 2.16 5.71 2.76 ;
        RECT  6.39 2.30 6.55 2.76 ;
        RECT  5.55 2.60 6.55 2.76 ;
    END
END HASP8V1_0

MACRO HASP4V1_0
    CLASS CORE ;
    FOREIGN HASP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.24 1.52 3.52 1.94 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.72 1.40 6.08 1.70 ;
        END
    END B
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 14.95  LAYER ME1  ;
        ANTENNADIFFAREA 7.28  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.71  LAYER ME1  ;
        ANTENNAMAXAREACAR 21.05  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.86 1.52 7.08 1.68 ;
        RECT  6.70 1.86 7.02 2.14 ;
        RECT  6.86 0.96 7.02 2.14 ;
        RECT  6.70 0.64 6.98 1.24 ;
        END
    END OUT
    PIN C
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 14.97  LAYER ME1  ;
        ANTENNADIFFAREA 7.29  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.71  LAYER ME1  ;
        ANTENNAMAXAREACAR 21.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.62 1.84 0.90 2.44 ;
        RECT  0.62 0.64 0.90 1.24 ;
        RECT  0.62 0.64 0.78 2.44 ;
        RECT  0.52 1.52 0.78 1.68 ;
        END
    END C
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 7.60 3.48 ;
        RECT  7.22 1.86 7.50 2.46 ;
        RECT  7.14 2.88 7.44 3.48 ;
        RECT  7.28 1.86 7.44 3.48 ;
        RECT  6.04 2.62 6.32 3.48 ;
        RECT  3.44 2.16 3.72 2.44 ;
        RECT  3.50 2.16 3.66 3.48 ;
        RECT  2.22 1.84 2.50 2.12 ;
        RECT  2.28 1.84 2.44 3.48 ;
        RECT  1.14 1.84 1.42 2.44 ;
        RECT  1.20 1.84 1.36 3.48 ;
        RECT  0.10 1.84 0.38 2.44 ;
        RECT  0.16 1.84 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 7.60 0.28 ;
        RECT  7.22 0.64 7.50 1.24 ;
        RECT  7.28 -0.28 7.44 1.24 ;
        RECT  7.14 -0.28 7.44 0.32 ;
        RECT  6.18 0.64 6.46 1.24 ;
        RECT  6.24 -0.28 6.40 1.24 ;
        RECT  3.16 0.76 3.44 1.04 ;
        RECT  3.22 -0.28 3.38 1.04 ;
        RECT  1.14 0.64 1.42 1.24 ;
        RECT  1.20 -0.28 1.36 1.24 ;
        RECT  0.10 0.64 0.38 1.24 ;
        RECT  0.16 -0.28 0.32 1.24 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  2.02 0.96 2.30 1.24 ;
        RECT  1.78 1.08 2.30 1.24 ;
        RECT  0.96 1.46 1.94 1.62 ;
        RECT  0.96 1.40 1.24 1.68 ;
        RECT  1.78 1.08 1.94 2.12 ;
        RECT  1.70 1.84 1.98 2.12 ;
        RECT  3.92 0.76 4.28 1.04 ;
        RECT  4.12 0.76 4.28 2.44 ;
        RECT  3.96 2.16 4.28 2.44 ;
        RECT  3.60 0.44 5.12 0.60 ;
        RECT  2.64 0.76 2.92 1.04 ;
        RECT  4.96 0.76 5.24 1.04 ;
        RECT  3.60 0.44 3.76 1.36 ;
        RECT  2.76 1.20 3.96 1.36 ;
        RECT  3.68 1.20 3.96 1.48 ;
        RECT  2.76 0.76 2.92 2.44 ;
        RECT  4.96 0.44 5.12 2.44 ;
        RECT  2.76 2.16 3.20 2.44 ;
        RECT  4.96 2.16 5.28 2.44 ;
        RECT  5.62 0.96 5.90 1.24 ;
        RECT  5.40 1.08 5.90 1.24 ;
        RECT  5.28 1.40 5.56 1.68 ;
        RECT  5.40 1.08 5.56 2.02 ;
        RECT  5.40 1.86 5.90 2.02 ;
        RECT  5.62 1.86 5.90 2.14 ;
        RECT  4.44 0.76 4.72 1.04 ;
        RECT  6.38 1.40 6.70 1.68 ;
        RECT  4.54 0.76 4.70 2.44 ;
        RECT  4.48 2.16 4.76 2.44 ;
        RECT  6.38 1.40 6.54 2.46 ;
        RECT  5.44 2.30 6.54 2.46 ;
        RECT  4.60 2.16 4.76 2.76 ;
        RECT  5.44 2.30 5.60 2.76 ;
        RECT  4.60 2.60 5.60 2.76 ;
    END
END HASP4V1_0

MACRO HASP2V1_0
    CLASS CORE ;
    FOREIGN HASP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN C
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 12.58  LAYER ME1  ;
        ANTENNADIFFAREA 5.70  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.42  LAYER ME1  ;
        ANTENNAMAXAREACAR 29.78  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.84 0.38 2.44 ;
        RECT  0.10 0.64 0.38 1.24 ;
        RECT  0.12 0.64 0.28 2.44 ;
        END
    END C
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 12.58  LAYER ME1  ;
        ANTENNADIFFAREA 5.70  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.42  LAYER ME1  ;
        ANTENNAMAXAREACAR 29.78  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.96 1.86 6.28 2.14 ;
        RECT  6.12 0.96 6.28 2.14 ;
        RECT  5.96 0.64 6.24 1.24 ;
        END
    END OUT
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.12 1.40 5.48 1.70 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.46 1.52 2.74 1.90 ;
        END
    END A
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 6.40 0.28 ;
        RECT  5.94 -0.28 6.22 0.32 ;
        RECT  5.44 0.64 5.72 1.24 ;
        RECT  5.50 -0.28 5.66 1.24 ;
        RECT  2.50 0.76 2.78 1.04 ;
        RECT  2.56 -0.28 2.72 1.04 ;
        RECT  0.62 0.64 0.90 1.24 ;
        RECT  0.68 -0.28 0.84 1.24 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 6.40 3.48 ;
        RECT  5.94 2.88 6.22 3.48 ;
        RECT  5.30 2.62 5.58 3.48 ;
        RECT  2.70 2.06 2.98 2.34 ;
        RECT  2.76 2.06 2.92 3.48 ;
        RECT  1.70 1.84 1.98 2.12 ;
        RECT  1.76 1.84 1.92 3.48 ;
        RECT  0.62 1.84 0.90 2.44 ;
        RECT  0.68 1.84 0.84 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  1.50 0.96 1.78 1.24 ;
        RECT  1.26 1.08 1.78 1.24 ;
        RECT  0.44 1.46 1.42 1.62 ;
        RECT  0.44 1.40 0.72 1.68 ;
        RECT  1.26 1.08 1.42 2.12 ;
        RECT  1.18 1.84 1.46 2.12 ;
        RECT  3.26 0.76 3.58 1.04 ;
        RECT  3.42 0.76 3.58 2.34 ;
        RECT  3.22 2.06 3.58 2.34 ;
        RECT  2.94 0.44 4.46 0.60 ;
        RECT  1.98 0.76 2.30 1.04 ;
        RECT  4.30 0.76 4.58 1.04 ;
        RECT  2.94 0.44 3.10 1.36 ;
        RECT  2.14 1.20 3.14 1.36 ;
        RECT  2.98 1.20 3.14 1.74 ;
        RECT  2.98 1.46 3.26 1.74 ;
        RECT  2.14 0.76 2.30 2.34 ;
        RECT  4.30 0.44 4.46 2.34 ;
        RECT  2.14 2.06 2.46 2.34 ;
        RECT  4.26 2.06 4.54 2.34 ;
        RECT  4.80 0.96 5.16 1.24 ;
        RECT  4.68 1.40 4.96 1.68 ;
        RECT  4.80 0.96 4.96 2.14 ;
        RECT  4.80 1.86 5.16 2.14 ;
        RECT  3.78 0.76 4.06 1.04 ;
        RECT  5.64 1.40 5.96 1.68 ;
        RECT  3.80 0.76 3.96 2.34 ;
        RECT  3.74 2.06 4.02 2.34 ;
        RECT  5.64 1.40 5.80 2.46 ;
        RECT  4.70 2.30 5.80 2.46 ;
        RECT  3.86 2.06 4.02 2.66 ;
        RECT  4.70 2.30 4.86 2.66 ;
        RECT  3.86 2.50 4.86 2.66 ;
    END
END HASP2V1_0

MACRO HASP1V1_0
    CLASS CORE ;
    FOREIGN HASP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.46 1.52 2.74 1.90 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.20 1.40 5.60 1.70 ;
        END
    END B
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 12.06  LAYER ME1  ;
        ANTENNADIFFAREA 4.85  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.27  LAYER ME1  ;
        ANTENNAMAXAREACAR 44.88  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.92 1.86 6.28 2.14 ;
        RECT  6.12 0.96 6.28 2.14 ;
        RECT  5.92 0.96 6.28 1.24 ;
        END
    END OUT
    PIN C
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 11.81  LAYER ME1  ;
        ANTENNADIFFAREA 4.96  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.27  LAYER ME1  ;
        ANTENNAMAXAREACAR 43.94  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.84 0.38 2.12 ;
        RECT  0.10 0.96 0.38 1.24 ;
        RECT  0.12 0.96 0.28 2.12 ;
        END
    END C
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 6.40 3.48 ;
        RECT  5.94 2.88 6.22 3.48 ;
        RECT  5.30 2.62 5.58 3.48 ;
        RECT  2.66 2.06 2.94 2.34 ;
        RECT  2.72 2.06 2.88 3.48 ;
        RECT  1.66 1.84 1.94 2.12 ;
        RECT  1.72 1.84 1.88 3.48 ;
        RECT  0.62 1.84 0.90 2.12 ;
        RECT  0.68 1.84 0.84 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 6.40 0.28 ;
        RECT  5.94 -0.28 6.22 0.32 ;
        RECT  5.40 0.96 5.68 1.24 ;
        RECT  5.46 -0.28 5.62 1.24 ;
        RECT  2.46 0.76 2.74 1.04 ;
        RECT  2.52 -0.28 2.68 1.04 ;
        RECT  0.62 0.96 0.90 1.24 ;
        RECT  0.68 -0.28 0.84 1.24 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  1.46 0.96 1.74 1.24 ;
        RECT  1.26 1.08 1.74 1.24 ;
        RECT  0.44 1.46 1.42 1.62 ;
        RECT  0.44 1.40 0.72 1.68 ;
        RECT  1.26 1.08 1.42 2.12 ;
        RECT  1.14 1.84 1.42 2.12 ;
        RECT  3.22 0.76 3.54 1.04 ;
        RECT  3.38 0.76 3.54 2.34 ;
        RECT  3.18 2.06 3.54 2.34 ;
        RECT  2.90 0.44 4.42 0.60 ;
        RECT  1.94 0.76 2.26 1.04 ;
        RECT  4.26 0.76 4.54 1.04 ;
        RECT  2.90 0.44 3.06 1.36 ;
        RECT  2.10 1.20 3.10 1.36 ;
        RECT  2.94 1.20 3.10 1.74 ;
        RECT  2.94 1.46 3.22 1.74 ;
        RECT  2.10 0.76 2.26 2.34 ;
        RECT  4.26 0.44 4.42 2.34 ;
        RECT  2.10 2.06 2.42 2.34 ;
        RECT  4.22 2.06 4.50 2.34 ;
        RECT  4.88 0.96 5.16 1.24 ;
        RECT  4.72 1.40 5.04 1.68 ;
        RECT  4.88 0.96 5.04 2.14 ;
        RECT  4.88 1.86 5.16 2.14 ;
        RECT  3.74 0.76 4.02 1.04 ;
        RECT  3.76 0.76 3.92 2.34 ;
        RECT  3.70 2.06 3.98 2.34 ;
        RECT  4.66 2.30 6.02 2.46 ;
        RECT  3.82 2.06 3.98 2.66 ;
        RECT  5.74 2.30 6.02 2.58 ;
        RECT  4.66 2.30 4.82 2.66 ;
        RECT  3.82 2.50 4.82 2.66 ;
    END
END HASP1V1_0

MACRO FILLER8EV1_0
    CLASS CORE ;
    FOREIGN FILLER8EV1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 3.20 3.48 ;
        RECT  2.72 2.88 3.02 3.48 ;
        RECT  2.72 1.86 3.00 3.48 ;
        RECT  2.12 1.86 2.40 3.48 ;
        RECT  1.52 1.86 1.80 3.48 ;
        RECT  0.92 1.86 1.20 3.48 ;
        RECT  0.22 1.86 0.60 2.14 ;
        RECT  0.22 1.38 0.50 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 3.20 0.28 ;
        RECT  2.82 -0.28 3.10 1.70 ;
        RECT  2.72 0.94 3.10 1.22 ;
        RECT  2.74 -0.28 3.10 0.32 ;
        RECT  2.12 -0.28 2.40 1.22 ;
        RECT  1.52 -0.28 1.80 1.22 ;
        RECT  0.92 -0.28 1.20 1.22 ;
        RECT  0.32 -0.28 0.60 1.22 ;
        END
    END GND!
END FILLER8EV1_0

MACRO FILLER64EV1_0
    CLASS CORE ;
    FOREIGN FILLER64EV1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 25.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 25.60 3.48 ;
        RECT  25.12 2.88 25.42 3.48 ;
        RECT  25.12 1.86 25.40 3.48 ;
        RECT  24.52 1.86 24.80 3.48 ;
        RECT  23.92 1.86 24.20 3.48 ;
        RECT  23.32 1.86 23.60 3.48 ;
        RECT  22.72 1.86 23.00 3.48 ;
        RECT  22.12 1.86 22.40 3.48 ;
        RECT  21.52 1.86 21.80 3.48 ;
        RECT  20.92 1.86 21.20 3.48 ;
        RECT  20.32 1.86 20.60 3.48 ;
        RECT  19.72 1.86 20.00 3.48 ;
        RECT  19.12 1.86 19.40 3.48 ;
        RECT  18.52 1.86 18.80 3.48 ;
        RECT  17.92 1.86 18.20 3.48 ;
        RECT  17.32 1.86 17.60 3.48 ;
        RECT  16.72 1.86 17.00 3.48 ;
        RECT  16.12 1.86 16.40 3.48 ;
        RECT  15.52 1.86 15.80 3.48 ;
        RECT  14.92 1.86 15.20 3.48 ;
        RECT  14.32 1.86 14.60 3.48 ;
        RECT  13.72 1.86 14.00 3.48 ;
        RECT  13.12 1.86 13.40 3.48 ;
        RECT  12.52 1.86 12.80 3.48 ;
        RECT  11.92 1.86 12.20 3.48 ;
        RECT  11.32 1.86 11.60 3.48 ;
        RECT  10.72 1.86 11.00 3.48 ;
        RECT  10.12 1.86 10.40 3.48 ;
        RECT  9.52 1.86 9.80 3.48 ;
        RECT  8.92 1.86 9.20 3.48 ;
        RECT  8.32 1.86 8.60 3.48 ;
        RECT  7.72 1.86 8.00 3.48 ;
        RECT  7.12 1.86 7.40 3.48 ;
        RECT  6.52 1.86 6.80 3.48 ;
        RECT  5.92 1.86 6.20 3.48 ;
        RECT  5.32 1.86 5.60 3.48 ;
        RECT  4.72 1.86 5.00 3.48 ;
        RECT  4.12 1.86 4.40 3.48 ;
        RECT  3.52 1.86 3.80 3.48 ;
        RECT  2.92 1.86 3.20 3.48 ;
        RECT  2.32 1.86 2.60 3.48 ;
        RECT  1.72 1.86 2.00 3.48 ;
        RECT  1.12 1.86 1.40 3.48 ;
        RECT  0.42 1.86 0.80 2.14 ;
        RECT  0.42 1.38 0.70 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 25.60 0.28 ;
        RECT  25.22 -0.28 25.50 1.70 ;
        RECT  25.12 0.94 25.50 1.22 ;
        RECT  25.14 -0.28 25.50 0.32 ;
        RECT  24.52 -0.28 24.80 1.22 ;
        RECT  23.92 -0.28 24.20 1.22 ;
        RECT  23.32 -0.28 23.60 1.22 ;
        RECT  22.72 -0.28 23.00 1.22 ;
        RECT  22.12 -0.28 22.40 1.22 ;
        RECT  21.52 -0.28 21.80 1.22 ;
        RECT  20.92 -0.28 21.20 1.22 ;
        RECT  20.32 -0.28 20.60 1.22 ;
        RECT  19.72 -0.28 20.00 1.22 ;
        RECT  19.12 -0.28 19.40 1.22 ;
        RECT  18.52 -0.28 18.80 1.22 ;
        RECT  17.92 -0.28 18.20 1.22 ;
        RECT  17.32 -0.28 17.60 1.22 ;
        RECT  16.72 -0.28 17.00 1.22 ;
        RECT  16.12 -0.28 16.40 1.22 ;
        RECT  15.52 -0.28 15.80 1.22 ;
        RECT  14.92 -0.28 15.20 1.22 ;
        RECT  14.32 -0.28 14.60 1.22 ;
        RECT  13.72 -0.28 14.00 1.22 ;
        RECT  13.12 -0.28 13.40 1.22 ;
        RECT  12.52 -0.28 12.80 1.22 ;
        RECT  11.92 -0.28 12.20 1.22 ;
        RECT  11.32 -0.28 11.60 1.22 ;
        RECT  10.72 -0.28 11.00 1.22 ;
        RECT  10.12 -0.28 10.40 1.22 ;
        RECT  9.52 -0.28 9.80 1.22 ;
        RECT  8.92 -0.28 9.20 1.22 ;
        RECT  8.32 -0.28 8.60 1.22 ;
        RECT  7.72 -0.28 8.00 1.22 ;
        RECT  7.12 -0.28 7.40 1.22 ;
        RECT  6.52 -0.28 6.80 1.22 ;
        RECT  5.92 -0.28 6.20 1.22 ;
        RECT  5.32 -0.28 5.60 1.22 ;
        RECT  4.72 -0.28 5.00 1.22 ;
        RECT  4.12 -0.28 4.40 1.22 ;
        RECT  3.52 -0.28 3.80 1.22 ;
        RECT  2.92 -0.28 3.20 1.22 ;
        RECT  2.32 -0.28 2.60 1.22 ;
        RECT  1.72 -0.28 2.00 1.22 ;
        RECT  1.12 -0.28 1.40 1.22 ;
        RECT  0.52 -0.28 0.80 1.22 ;
        END
    END GND!
END FILLER64EV1_0

MACRO FILLER4EV1_0
    CLASS CORE ;
    FOREIGN FILLER4EV1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 1.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 1.60 3.48 ;
        RECT  1.16 2.26 1.44 2.54 ;
        RECT  1.14 2.88 1.42 3.48 ;
        RECT  1.22 2.26 1.38 3.48 ;
        RECT  0.56 1.54 0.84 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 1.60 0.28 ;
        RECT  1.16 0.66 1.44 1.82 ;
        RECT  1.14 -0.28 1.42 0.32 ;
        RECT  1.22 -0.28 1.38 1.82 ;
        RECT  0.56 -0.28 0.84 0.94 ;
        END
    END GND!
END FILLER4EV1_0

MACRO FILLER3V1_0
    CLASS CORE ;
    FOREIGN FILLER3V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 1.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 1.20 3.48 ;
        RECT  0.74 2.88 1.02 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 1.20 0.28 ;
        RECT  0.74 -0.28 1.02 0.32 ;
        END
    END GND!
END FILLER3V1_0

MACRO FILLER32EV1_0
    CLASS CORE ;
    FOREIGN FILLER32EV1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 12.80 0.28 ;
        RECT  12.42 -0.28 12.70 1.70 ;
        RECT  12.32 0.94 12.70 1.22 ;
        RECT  12.34 -0.28 12.70 0.32 ;
        RECT  11.72 -0.28 12.00 1.22 ;
        RECT  11.12 -0.28 11.40 1.22 ;
        RECT  10.52 -0.28 10.80 1.22 ;
        RECT  9.92 -0.28 10.20 1.22 ;
        RECT  9.32 -0.28 9.60 1.22 ;
        RECT  8.72 -0.28 9.00 1.22 ;
        RECT  8.12 -0.28 8.40 1.22 ;
        RECT  7.52 -0.28 7.80 1.22 ;
        RECT  6.92 -0.28 7.20 1.22 ;
        RECT  6.32 -0.28 6.60 1.22 ;
        RECT  5.72 -0.28 6.00 1.22 ;
        RECT  5.12 -0.28 5.40 1.22 ;
        RECT  4.52 -0.28 4.80 1.22 ;
        RECT  3.92 -0.28 4.20 1.22 ;
        RECT  3.32 -0.28 3.60 1.22 ;
        RECT  2.72 -0.28 3.00 1.22 ;
        RECT  2.12 -0.28 2.40 1.22 ;
        RECT  1.52 -0.28 1.80 1.22 ;
        RECT  0.92 -0.28 1.20 1.22 ;
        RECT  0.32 -0.28 0.60 1.22 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 12.80 3.48 ;
        RECT  12.32 2.88 12.62 3.48 ;
        RECT  12.32 1.86 12.60 3.48 ;
        RECT  11.72 1.86 12.00 3.48 ;
        RECT  11.12 1.86 11.40 3.48 ;
        RECT  10.52 1.86 10.80 3.48 ;
        RECT  9.92 1.86 10.20 3.48 ;
        RECT  9.32 1.86 9.60 3.48 ;
        RECT  8.72 1.86 9.00 3.48 ;
        RECT  8.12 1.86 8.40 3.48 ;
        RECT  7.52 1.86 7.80 3.48 ;
        RECT  6.92 1.86 7.20 3.48 ;
        RECT  6.32 1.86 6.60 3.48 ;
        RECT  5.72 1.86 6.00 3.48 ;
        RECT  5.12 1.86 5.40 3.48 ;
        RECT  4.52 1.86 4.80 3.48 ;
        RECT  3.92 1.86 4.20 3.48 ;
        RECT  3.32 1.86 3.60 3.48 ;
        RECT  2.72 1.86 3.00 3.48 ;
        RECT  2.12 1.86 2.40 3.48 ;
        RECT  1.52 1.86 1.80 3.48 ;
        RECT  0.92 1.86 1.20 3.48 ;
        RECT  0.22 1.86 0.60 2.14 ;
        RECT  0.22 1.38 0.50 3.48 ;
        END
    END VDD!
END FILLER32EV1_0

MACRO FILLER2V1_0
    CLASS CORE ;
    FOREIGN FILLER2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 0.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 0.80 3.48 ;
        RECT  0.34 2.88 0.62 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 0.80 0.28 ;
        RECT  0.34 -0.28 0.62 0.32 ;
        END
    END GND!
END FILLER2V1_0

MACRO FILLER1V1_0
    CLASS CORE ;
    FOREIGN FILLER1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 0.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 0.40 0.28 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 0.40 3.48 ;
        END
    END VDD!
END FILLER1V1_0

MACRO FILLER16EV1_0
    CLASS CORE ;
    FOREIGN FILLER16EV1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 6.40 3.48 ;
        RECT  5.92 2.88 6.22 3.48 ;
        RECT  5.92 1.86 6.20 3.48 ;
        RECT  5.32 1.86 5.60 3.48 ;
        RECT  4.72 1.86 5.00 3.48 ;
        RECT  4.12 1.86 4.40 3.48 ;
        RECT  3.52 1.86 3.80 3.48 ;
        RECT  2.92 1.86 3.20 3.48 ;
        RECT  2.32 1.86 2.60 3.48 ;
        RECT  1.72 1.86 2.00 3.48 ;
        RECT  1.12 1.86 1.40 3.48 ;
        RECT  0.42 1.86 0.80 2.14 ;
        RECT  0.42 1.38 0.70 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 6.40 0.28 ;
        RECT  6.02 -0.28 6.30 1.70 ;
        RECT  5.92 0.94 6.30 1.22 ;
        RECT  5.94 -0.28 6.30 0.32 ;
        RECT  5.32 -0.28 5.60 1.22 ;
        RECT  4.72 -0.28 5.00 1.22 ;
        RECT  4.12 -0.28 4.40 1.22 ;
        RECT  3.52 -0.28 3.80 1.22 ;
        RECT  2.92 -0.28 3.20 1.22 ;
        RECT  2.32 -0.28 2.60 1.22 ;
        RECT  1.72 -0.28 2.00 1.22 ;
        RECT  1.12 -0.28 1.40 1.22 ;
        RECT  0.52 -0.28 0.80 1.22 ;
        END
    END GND!
END FILLER16EV1_0

MACRO FASP8V1_0
    CLASS CORE ;
    FOREIGN FASP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 13.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 26.33  LAYER ME1  ;
        ANTENNADIFFAREA 13.35  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.56  LAYER ME1  ;
        ANTENNAMAXAREACAR 16.93  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.98 1.92 12.26 2.52 ;
        RECT  11.98 0.64 12.26 1.24 ;
        RECT  11.98 0.64 12.14 2.52 ;
        RECT  11.06 1.52 12.14 1.68 ;
        RECT  11.06 1.46 11.54 1.74 ;
        RECT  10.94 1.92 11.22 2.52 ;
        RECT  11.06 0.64 11.22 2.52 ;
        RECT  10.94 0.64 11.22 1.24 ;
        END
    END OUT
    PIN CI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.28 1.46 10.70 1.74 ;
        END
    END CI
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.27  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.50 1.46 7.92 1.74 ;
        END
    END B
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 26.33  LAYER ME1  ;
        ANTENNADIFFAREA 12.87  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.56  LAYER ME1  ;
        ANTENNAMAXAREACAR 16.93  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.66 1.96 1.94 2.56 ;
        RECT  1.66 0.56 1.94 1.16 ;
        RECT  1.66 0.56 1.82 2.56 ;
        RECT  0.68 1.52 1.82 1.68 ;
        RECT  0.68 1.46 1.14 1.74 ;
        RECT  0.62 1.96 0.90 2.56 ;
        RECT  0.62 0.56 0.90 1.16 ;
        RECT  0.68 0.56 0.84 2.56 ;
        END
    END CO
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 26.33  LAYER ME1  ;
        ANTENNADIFFAREA 12.73  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.56  LAYER ME1  ;
        ANTENNAMAXAREACAR 16.93  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.72 1.92 7.00 2.20 ;
        RECT  6.72 0.76 7.00 1.04 ;
        RECT  6.72 0.44 6.88 2.20 ;
        RECT  5.36 0.44 6.88 0.60 ;
        RECT  5.10 1.46 5.52 1.74 ;
        RECT  5.36 0.44 5.52 1.74 ;
        END
    END A
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 13.20 0.28 ;
        RECT  12.58 -0.28 13.02 0.32 ;
        RECT  12.50 0.64 12.78 1.24 ;
        RECT  12.58 -0.28 12.74 1.24 ;
        RECT  11.46 0.64 11.74 1.24 ;
        RECT  11.52 -0.28 11.68 1.24 ;
        RECT  10.42 0.64 10.70 1.24 ;
        RECT  10.48 -0.28 10.64 1.24 ;
        RECT  7.72 0.76 8.00 1.04 ;
        RECT  7.78 -0.28 7.94 1.04 ;
        RECT  4.92 -0.28 5.20 0.68 ;
        RECT  4.16 0.88 4.44 1.16 ;
        RECT  4.22 -0.28 4.38 1.16 ;
        RECT  2.18 0.56 2.46 1.16 ;
        RECT  2.24 -0.28 2.40 1.16 ;
        RECT  1.14 0.56 1.42 1.16 ;
        RECT  1.20 -0.28 1.36 1.16 ;
        RECT  0.10 0.56 0.38 1.16 ;
        RECT  0.16 -0.28 0.32 1.16 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 13.20 3.48 ;
        RECT  12.58 2.88 13.02 3.48 ;
        RECT  12.50 1.92 12.78 2.52 ;
        RECT  12.58 1.92 12.74 3.48 ;
        RECT  11.46 1.92 11.74 2.52 ;
        RECT  11.52 1.92 11.68 3.48 ;
        RECT  10.42 1.92 10.70 2.52 ;
        RECT  10.48 1.92 10.64 3.48 ;
        RECT  7.72 1.92 8.00 2.20 ;
        RECT  7.74 1.92 7.90 3.48 ;
        RECT  5.16 1.92 5.44 2.20 ;
        RECT  5.22 1.92 5.38 3.48 ;
        RECT  4.16 1.96 4.44 2.24 ;
        RECT  4.22 1.96 4.38 3.48 ;
        RECT  2.18 1.96 2.46 2.56 ;
        RECT  2.24 1.96 2.40 3.48 ;
        RECT  1.14 1.96 1.42 2.56 ;
        RECT  1.20 1.96 1.36 3.48 ;
        RECT  0.10 1.96 0.38 2.56 ;
        RECT  0.16 1.96 0.32 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  3.26 0.88 3.54 1.16 ;
        RECT  2.04 1.48 3.48 1.64 ;
        RECT  2.04 1.42 2.32 1.70 ;
        RECT  3.32 0.88 3.48 2.24 ;
        RECT  3.26 1.96 3.54 2.24 ;
        RECT  3.70 1.64 4.84 1.80 ;
        RECT  4.68 1.64 4.84 2.24 ;
        RECT  2.74 1.96 3.02 2.24 ;
        RECT  4.68 1.96 4.96 2.24 ;
        RECT  2.86 1.96 3.02 2.56 ;
        RECT  3.70 1.64 3.86 2.56 ;
        RECT  2.86 2.40 3.86 2.56 ;
        RECT  2.86 0.56 3.86 0.72 ;
        RECT  2.86 0.56 3.02 1.16 ;
        RECT  2.74 0.88 3.02 1.16 ;
        RECT  4.68 0.88 4.96 1.16 ;
        RECT  3.70 0.56 3.86 1.48 ;
        RECT  4.68 0.88 4.84 1.48 ;
        RECT  3.70 1.32 4.84 1.48 ;
        RECT  5.68 0.76 5.96 1.04 ;
        RECT  5.80 0.76 5.96 2.20 ;
        RECT  5.68 1.92 5.96 2.20 ;
        RECT  6.20 0.76 6.48 1.04 ;
        RECT  6.20 1.92 6.48 2.20 ;
        RECT  6.26 0.76 6.42 2.58 ;
        RECT  6.26 2.42 7.24 2.58 ;
        RECT  6.96 2.42 7.24 2.70 ;
        RECT  7.18 0.76 7.48 1.04 ;
        RECT  7.06 1.22 7.34 1.50 ;
        RECT  7.18 0.76 7.34 2.20 ;
        RECT  7.18 1.92 7.48 2.20 ;
        RECT  8.24 0.76 8.52 1.04 ;
        RECT  8.30 0.76 8.46 2.20 ;
        RECT  8.24 1.92 8.52 2.20 ;
        RECT  9.26 0.76 9.56 1.04 ;
        RECT  9.26 1.92 9.56 2.20 ;
        RECT  9.26 0.76 9.42 2.58 ;
        RECT  8.06 2.42 9.42 2.58 ;
        RECT  8.06 2.42 8.34 2.70 ;
        RECT  8.88 0.44 10.00 0.60 ;
        RECT  9.72 0.44 10.00 0.72 ;
        RECT  8.88 0.44 9.04 1.04 ;
        RECT  8.76 0.76 9.04 1.04 ;
        RECT  8.82 0.76 8.98 2.20 ;
        RECT  8.76 1.92 9.04 2.20 ;
        RECT  9.74 0.96 10.14 1.24 ;
        RECT  9.74 1.92 10.14 2.20 ;
        RECT  9.74 0.96 9.90 2.70 ;
        RECT  9.68 2.42 9.96 2.70 ;
    END
END FASP8V1_0

MACRO FASP4V1_0
    CLASS CORE ;
    FOREIGN FASP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 21.59  LAYER ME1  ;
        ANTENNADIFFAREA 10.18  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.98  LAYER ME1  ;
        ANTENNAMAXAREACAR 22.05  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.02 1.46 10.34 1.74 ;
        RECT  9.90 1.92 10.18 2.52 ;
        RECT  10.02 0.64 10.18 2.52 ;
        RECT  9.90 0.64 10.18 1.24 ;
        END
    END OUT
    PIN CI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.24 1.46 9.66 1.74 ;
        END
    END CI
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.27  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.46 1.46 6.88 1.74 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 21.59  LAYER ME1  ;
        ANTENNADIFFAREA 10.04  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.98  LAYER ME1  ;
        ANTENNAMAXAREACAR 22.05  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.68 1.92 5.96 2.20 ;
        RECT  5.68 0.76 5.96 1.04 ;
        RECT  5.68 0.44 5.84 2.20 ;
        RECT  4.32 0.44 5.84 0.60 ;
        RECT  4.06 1.46 4.48 1.74 ;
        RECT  4.32 0.44 4.48 1.74 ;
        END
    END A
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 21.59  LAYER ME1  ;
        ANTENNADIFFAREA 9.71  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.98  LAYER ME1  ;
        ANTENNAMAXAREACAR 22.05  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.62 1.96 0.90 2.56 ;
        RECT  0.62 0.56 0.90 1.16 ;
        RECT  0.62 0.56 0.78 2.56 ;
        RECT  0.46 1.46 0.78 1.74 ;
        END
    END CO
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 10.80 0.28 ;
        RECT  10.42 0.64 10.70 1.24 ;
        RECT  10.48 -0.28 10.64 1.24 ;
        RECT  10.34 -0.28 10.64 0.32 ;
        RECT  9.38 0.64 9.66 1.24 ;
        RECT  9.44 -0.28 9.60 1.24 ;
        RECT  6.68 0.76 6.96 1.04 ;
        RECT  6.74 -0.28 6.90 1.04 ;
        RECT  3.88 -0.28 4.16 0.68 ;
        RECT  3.12 0.88 3.40 1.16 ;
        RECT  3.18 -0.28 3.34 1.16 ;
        RECT  1.14 0.56 1.42 1.16 ;
        RECT  1.20 -0.28 1.36 1.16 ;
        RECT  0.10 0.56 0.38 1.16 ;
        RECT  0.16 -0.28 0.32 1.16 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 10.80 3.48 ;
        RECT  10.42 1.92 10.70 2.52 ;
        RECT  10.34 2.88 10.64 3.48 ;
        RECT  10.48 1.92 10.64 3.48 ;
        RECT  9.38 1.92 9.66 2.52 ;
        RECT  9.44 1.92 9.60 3.48 ;
        RECT  6.68 1.92 6.96 2.20 ;
        RECT  6.70 1.92 6.86 3.48 ;
        RECT  4.12 1.92 4.40 2.20 ;
        RECT  4.18 1.92 4.34 3.48 ;
        RECT  3.12 1.96 3.40 2.24 ;
        RECT  3.18 1.96 3.34 3.48 ;
        RECT  1.14 1.96 1.42 2.56 ;
        RECT  1.20 1.96 1.36 3.48 ;
        RECT  0.10 1.96 0.38 2.56 ;
        RECT  0.16 1.96 0.32 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  2.22 0.88 2.50 1.16 ;
        RECT  1.00 1.48 2.44 1.64 ;
        RECT  1.00 1.42 1.28 1.70 ;
        RECT  2.28 0.88 2.44 2.24 ;
        RECT  2.22 1.96 2.50 2.24 ;
        RECT  2.66 1.64 3.80 1.80 ;
        RECT  3.64 1.64 3.80 2.24 ;
        RECT  1.70 1.96 1.98 2.24 ;
        RECT  3.64 1.96 3.92 2.24 ;
        RECT  1.82 1.96 1.98 2.56 ;
        RECT  2.66 1.64 2.82 2.56 ;
        RECT  1.82 2.40 2.82 2.56 ;
        RECT  1.82 0.56 2.82 0.72 ;
        RECT  1.82 0.56 1.98 1.16 ;
        RECT  1.70 0.88 1.98 1.16 ;
        RECT  3.64 0.88 3.92 1.16 ;
        RECT  2.66 0.56 2.82 1.48 ;
        RECT  3.64 0.88 3.80 1.48 ;
        RECT  2.66 1.32 3.80 1.48 ;
        RECT  4.64 0.76 4.92 1.04 ;
        RECT  4.76 0.76 4.92 2.20 ;
        RECT  4.64 1.92 4.92 2.20 ;
        RECT  5.16 0.76 5.44 1.04 ;
        RECT  5.16 1.92 5.44 2.20 ;
        RECT  5.22 0.76 5.38 2.58 ;
        RECT  5.22 2.42 6.20 2.58 ;
        RECT  5.92 2.42 6.20 2.70 ;
        RECT  6.14 0.76 6.44 1.04 ;
        RECT  6.02 1.22 6.30 1.50 ;
        RECT  6.14 0.76 6.30 2.20 ;
        RECT  6.14 1.92 6.44 2.20 ;
        RECT  7.20 0.76 7.48 1.04 ;
        RECT  7.26 0.76 7.42 2.20 ;
        RECT  7.20 1.92 7.48 2.20 ;
        RECT  8.22 0.76 8.52 1.04 ;
        RECT  8.22 1.92 8.52 2.20 ;
        RECT  8.22 0.76 8.38 2.58 ;
        RECT  7.02 2.42 8.38 2.58 ;
        RECT  7.02 2.42 7.30 2.70 ;
        RECT  7.84 0.44 8.96 0.60 ;
        RECT  8.68 0.44 8.96 0.72 ;
        RECT  7.84 0.44 8.00 1.04 ;
        RECT  7.72 0.76 8.00 1.04 ;
        RECT  7.78 0.76 7.94 2.20 ;
        RECT  7.72 1.92 8.00 2.20 ;
        RECT  8.70 0.96 9.10 1.24 ;
        RECT  8.70 1.92 9.10 2.20 ;
        RECT  8.70 0.96 8.86 2.70 ;
        RECT  8.64 2.42 8.92 2.70 ;
    END
END FASP4V1_0

MACRO FASP2V1_0
    CLASS CORE ;
    FOREIGN FASP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 19.77  LAYER ME1  ;
        ANTENNADIFFAREA 8.69  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.69  LAYER ME1  ;
        ANTENNAMAXAREACAR 28.60  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.50 1.46 9.92 1.74 ;
        RECT  9.38 1.92 9.66 2.52 ;
        RECT  9.50 0.64 9.66 2.52 ;
        RECT  9.38 0.64 9.66 1.24 ;
        END
    END OUT
    PIN CI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.72 1.46 9.14 1.74 ;
        END
    END CI
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 19.77  LAYER ME1  ;
        ANTENNADIFFAREA 8.79  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.69  LAYER ME1  ;
        ANTENNAMAXAREACAR 28.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.16 1.92 5.44 2.20 ;
        RECT  5.16 0.76 5.44 1.04 ;
        RECT  5.16 0.44 5.32 2.20 ;
        RECT  3.80 0.44 5.32 0.60 ;
        RECT  3.66 1.40 3.96 1.76 ;
        RECT  3.80 0.44 3.96 1.76 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.27  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.98 1.46 6.38 1.74 ;
        END
    END B
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 19.77  LAYER ME1  ;
        ANTENNADIFFAREA 8.49  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.69  LAYER ME1  ;
        ANTENNAMAXAREACAR 28.60  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.96 0.38 2.56 ;
        RECT  0.10 0.56 0.38 1.16 ;
        RECT  0.12 0.56 0.28 2.56 ;
        END
    END CO
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 10.00 3.48 ;
        RECT  9.54 2.88 9.82 3.48 ;
        RECT  8.86 1.92 9.14 2.52 ;
        RECT  8.92 1.92 9.08 3.48 ;
        RECT  6.16 1.92 6.44 2.20 ;
        RECT  6.18 1.92 6.34 3.48 ;
        RECT  3.60 1.92 3.88 2.20 ;
        RECT  3.66 1.92 3.82 3.48 ;
        RECT  2.60 1.96 2.88 2.24 ;
        RECT  2.66 1.96 2.82 3.48 ;
        RECT  0.62 1.96 0.90 2.56 ;
        RECT  0.68 1.96 0.84 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 10.00 0.28 ;
        RECT  9.54 -0.28 9.82 0.32 ;
        RECT  8.86 0.64 9.14 1.24 ;
        RECT  8.92 -0.28 9.08 1.24 ;
        RECT  6.16 0.76 6.44 1.04 ;
        RECT  6.22 -0.28 6.38 1.04 ;
        RECT  3.36 -0.28 3.64 0.68 ;
        RECT  2.60 0.88 2.88 1.16 ;
        RECT  2.66 -0.28 2.82 1.16 ;
        RECT  0.62 0.56 0.90 1.16 ;
        RECT  0.68 -0.28 0.84 1.16 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  1.70 0.88 1.98 1.16 ;
        RECT  0.48 1.48 1.92 1.64 ;
        RECT  0.48 1.42 0.76 1.70 ;
        RECT  1.76 0.88 1.92 2.24 ;
        RECT  1.70 1.96 1.98 2.24 ;
        RECT  2.14 1.64 3.28 1.80 ;
        RECT  3.12 1.64 3.28 2.24 ;
        RECT  1.18 1.96 1.46 2.24 ;
        RECT  3.12 1.96 3.40 2.24 ;
        RECT  1.30 1.96 1.46 2.56 ;
        RECT  2.14 1.64 2.30 2.56 ;
        RECT  1.30 2.40 2.30 2.56 ;
        RECT  1.30 0.56 2.30 0.72 ;
        RECT  1.30 0.56 1.46 1.16 ;
        RECT  1.18 0.88 1.46 1.16 ;
        RECT  3.12 0.88 3.40 1.16 ;
        RECT  2.14 0.56 2.30 1.48 ;
        RECT  3.12 0.88 3.28 1.48 ;
        RECT  2.14 1.32 3.28 1.48 ;
        RECT  4.12 0.76 4.40 1.04 ;
        RECT  4.24 0.76 4.40 2.20 ;
        RECT  4.12 1.92 4.40 2.20 ;
        RECT  4.64 0.76 4.92 1.04 ;
        RECT  4.64 1.92 4.92 2.20 ;
        RECT  4.70 0.76 4.86 2.58 ;
        RECT  4.70 2.42 5.68 2.58 ;
        RECT  5.40 2.42 5.68 2.70 ;
        RECT  5.64 0.76 5.92 1.04 ;
        RECT  5.50 1.22 5.80 1.50 ;
        RECT  5.64 0.76 5.80 2.20 ;
        RECT  5.64 1.92 5.92 2.20 ;
        RECT  6.68 0.76 6.96 1.04 ;
        RECT  6.74 0.76 6.90 2.20 ;
        RECT  6.68 1.92 6.96 2.20 ;
        RECT  7.70 0.76 8.00 1.04 ;
        RECT  7.70 1.92 8.00 2.20 ;
        RECT  7.70 0.76 7.86 2.58 ;
        RECT  6.50 2.42 7.86 2.58 ;
        RECT  6.50 2.42 6.78 2.70 ;
        RECT  7.32 0.44 8.44 0.60 ;
        RECT  8.16 0.44 8.44 0.72 ;
        RECT  7.32 0.44 7.48 1.04 ;
        RECT  7.20 0.76 7.48 1.04 ;
        RECT  7.26 0.76 7.42 2.20 ;
        RECT  7.20 1.92 7.48 2.20 ;
        RECT  8.18 0.96 8.58 1.24 ;
        RECT  8.18 1.92 8.58 2.20 ;
        RECT  8.18 0.96 8.34 2.70 ;
        RECT  8.12 2.42 8.40 2.70 ;
    END
END FASP2V1_0

MACRO FASP1V1_0
    CLASS CORE ;
    FOREIGN FASP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 19.24  LAYER ME1  ;
        ANTENNADIFFAREA 7.69  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.54  LAYER ME1  ;
        ANTENNAMAXAREACAR 35.79  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.30 1.92 9.58 2.20 ;
        RECT  9.30 0.96 9.58 1.24 ;
        RECT  9.30 0.96 9.54 2.20 ;
        RECT  9.26 1.46 9.54 1.74 ;
        END
    END OUT
    PIN CI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.46 1.40 8.78 1.76 ;
        END
    END CI
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 18.96  LAYER ME1  ;
        ANTENNADIFFAREA 7.58  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.54  LAYER ME1  ;
        ANTENNAMAXAREACAR 35.26  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.96 0.38 2.24 ;
        RECT  0.10 0.88 0.38 1.16 ;
        RECT  0.12 0.88 0.28 2.24 ;
        END
    END CO
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.27  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.94 1.46 6.34 1.74 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 19.24  LAYER ME1  ;
        ANTENNADIFFAREA 7.78  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.54  LAYER ME1  ;
        ANTENNAMAXAREACAR 35.79  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.12 1.92 5.40 2.20 ;
        RECT  5.12 0.76 5.40 1.04 ;
        RECT  5.12 0.44 5.28 2.20 ;
        RECT  3.76 0.44 5.28 0.60 ;
        RECT  3.66 1.40 3.94 1.76 ;
        RECT  3.76 0.44 3.92 1.76 ;
        END
    END A
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 10.00 0.28 ;
        RECT  9.54 -0.28 9.82 0.32 ;
        RECT  8.78 0.96 9.06 1.24 ;
        RECT  8.84 -0.28 9.00 1.24 ;
        RECT  6.12 0.76 6.40 1.04 ;
        RECT  6.18 -0.28 6.34 1.04 ;
        RECT  3.32 -0.28 3.60 0.68 ;
        RECT  2.56 0.88 2.84 1.16 ;
        RECT  2.62 -0.28 2.78 1.16 ;
        RECT  0.62 0.88 0.90 1.16 ;
        RECT  0.68 -0.28 0.84 1.16 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 10.00 3.48 ;
        RECT  9.54 2.88 9.82 3.48 ;
        RECT  8.78 1.92 9.06 2.20 ;
        RECT  8.84 1.92 9.00 3.48 ;
        RECT  6.12 1.92 6.40 2.20 ;
        RECT  6.14 1.92 6.30 3.48 ;
        RECT  3.56 1.92 3.84 2.20 ;
        RECT  3.62 1.92 3.78 3.48 ;
        RECT  2.56 1.96 2.84 2.24 ;
        RECT  2.62 1.96 2.78 3.48 ;
        RECT  0.62 1.96 0.90 2.24 ;
        RECT  0.68 1.96 0.84 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  1.66 0.88 1.94 1.16 ;
        RECT  0.44 1.48 1.88 1.64 ;
        RECT  0.44 1.42 0.72 1.70 ;
        RECT  1.72 0.88 1.88 2.24 ;
        RECT  1.66 1.96 1.94 2.24 ;
        RECT  2.10 1.64 3.24 1.80 ;
        RECT  3.08 1.64 3.24 2.24 ;
        RECT  1.14 1.96 1.42 2.24 ;
        RECT  3.08 1.96 3.36 2.24 ;
        RECT  1.26 1.96 1.42 2.56 ;
        RECT  2.10 1.64 2.26 2.56 ;
        RECT  1.26 2.40 2.26 2.56 ;
        RECT  1.26 0.56 2.26 0.72 ;
        RECT  1.26 0.56 1.42 1.16 ;
        RECT  1.14 0.88 1.42 1.16 ;
        RECT  3.08 0.88 3.36 1.16 ;
        RECT  2.10 0.56 2.26 1.48 ;
        RECT  3.08 0.88 3.24 1.48 ;
        RECT  2.10 1.32 3.24 1.48 ;
        RECT  4.08 0.76 4.36 1.04 ;
        RECT  4.20 0.76 4.36 2.20 ;
        RECT  4.08 1.92 4.36 2.20 ;
        RECT  4.60 0.76 4.88 1.04 ;
        RECT  4.60 1.92 4.88 2.20 ;
        RECT  4.66 0.76 4.82 2.58 ;
        RECT  4.66 2.42 5.64 2.58 ;
        RECT  5.36 2.42 5.64 2.70 ;
        RECT  5.60 0.76 5.88 1.04 ;
        RECT  5.46 1.22 5.76 1.50 ;
        RECT  5.60 0.76 5.76 2.20 ;
        RECT  5.60 1.92 5.88 2.20 ;
        RECT  6.64 0.76 6.92 1.04 ;
        RECT  6.70 0.76 6.86 2.20 ;
        RECT  6.64 1.92 6.92 2.20 ;
        RECT  7.66 0.76 7.96 1.04 ;
        RECT  7.66 1.92 7.96 2.20 ;
        RECT  7.66 0.76 7.82 2.58 ;
        RECT  6.46 2.42 7.82 2.58 ;
        RECT  6.46 2.42 6.74 2.70 ;
        RECT  7.28 0.44 8.40 0.60 ;
        RECT  8.12 0.44 8.40 0.72 ;
        RECT  7.28 0.44 7.44 1.04 ;
        RECT  7.16 0.76 7.44 1.04 ;
        RECT  7.22 0.76 7.38 2.20 ;
        RECT  7.16 1.92 7.44 2.20 ;
        RECT  8.14 0.96 8.54 1.24 ;
        RECT  8.14 1.92 8.54 2.20 ;
        RECT  8.14 0.96 8.30 2.70 ;
        RECT  8.08 2.42 8.36 2.70 ;
    END
END FASP1V1_0

MACRO DLAHSP8V1_0
    CLASS CORE ;
    FOREIGN DLAHSP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 19.33  LAYER ME1  ;
        ANTENNADIFFAREA 10.12  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.60  LAYER ME1  ;
        ANTENNAMAXAREACAR 12.06  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.88 1.84 9.16 2.50 ;
        RECT  8.88 0.58 9.16 1.24 ;
        RECT  8.92 0.58 9.08 2.50 ;
        RECT  7.96 1.52 9.08 1.68 ;
        RECT  7.84 1.84 8.12 2.50 ;
        RECT  7.96 0.58 8.12 2.50 ;
        RECT  7.84 0.58 8.12 1.24 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 19.33  LAYER ME1  ;
        ANTENNADIFFAREA 10.92  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.60  LAYER ME1  ;
        ANTENNAMAXAREACAR 12.06  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.80 1.84 7.08 2.50 ;
        RECT  6.80 0.58 7.08 1.24 ;
        RECT  6.80 0.58 6.96 2.50 ;
        RECT  5.72 1.52 6.96 1.68 ;
        RECT  5.72 1.84 6.04 2.50 ;
        RECT  5.72 0.58 6.04 1.24 ;
        RECT  5.72 0.58 5.88 2.50 ;
        END
    END QB
    PIN G
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.32 1.40 0.74 1.68 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.99 1.46 2.41 1.74 ;
        END
    END D
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 10.00 0.28 ;
        RECT  9.46 -0.28 9.82 0.32 ;
        RECT  9.40 0.58 9.68 1.24 ;
        RECT  9.46 -0.28 9.62 1.24 ;
        RECT  8.36 0.58 8.64 1.24 ;
        RECT  8.42 -0.28 8.58 1.24 ;
        RECT  7.32 0.58 7.60 1.24 ;
        RECT  7.38 -0.28 7.54 1.24 ;
        RECT  6.28 0.58 6.56 1.24 ;
        RECT  6.34 -0.28 6.50 1.24 ;
        RECT  5.24 0.58 5.52 1.24 ;
        RECT  5.30 -0.28 5.46 1.24 ;
        RECT  4.24 0.73 4.52 1.01 ;
        RECT  4.30 -0.28 4.46 1.01 ;
        RECT  1.92 0.73 2.20 1.01 ;
        RECT  1.98 -0.28 2.14 1.01 ;
        RECT  0.22 0.96 0.50 1.24 ;
        RECT  0.28 -0.28 0.44 1.24 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 10.00 3.48 ;
        RECT  9.46 2.88 9.82 3.48 ;
        RECT  9.40 1.84 9.68 2.50 ;
        RECT  9.46 1.84 9.62 3.48 ;
        RECT  8.36 1.84 8.64 2.50 ;
        RECT  8.42 1.84 8.58 3.48 ;
        RECT  7.32 1.84 7.60 2.50 ;
        RECT  7.38 1.84 7.54 3.48 ;
        RECT  6.28 1.84 6.56 2.50 ;
        RECT  6.34 1.84 6.50 3.48 ;
        RECT  5.24 1.84 5.52 2.50 ;
        RECT  5.30 1.84 5.46 3.48 ;
        RECT  4.24 1.90 4.52 2.18 ;
        RECT  4.30 1.90 4.46 3.48 ;
        RECT  1.92 1.90 2.20 2.18 ;
        RECT  1.98 1.90 2.14 3.48 ;
        RECT  0.22 1.84 0.50 2.12 ;
        RECT  0.29 1.84 0.45 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.74 0.96 1.06 1.24 ;
        RECT  0.90 1.40 1.30 1.68 ;
        RECT  0.90 0.96 1.06 2.12 ;
        RECT  0.74 1.84 1.06 2.12 ;
        RECT  1.40 0.73 1.68 1.01 ;
        RECT  1.46 0.73 1.62 2.18 ;
        RECT  1.34 1.90 1.68 2.18 ;
        RECT  1.34 1.90 1.50 2.76 ;
        RECT  1.22 2.48 1.50 2.76 ;
        RECT  2.44 0.73 2.77 1.01 ;
        RECT  2.61 0.73 2.77 2.18 ;
        RECT  2.44 1.90 2.77 2.18 ;
        RECT  3.48 0.73 3.76 1.01 ;
        RECT  3.54 0.73 3.70 2.18 ;
        RECT  3.48 1.90 3.76 2.18 ;
        RECT  2.96 0.73 3.24 1.01 ;
        RECT  2.96 1.90 3.24 2.18 ;
        RECT  3.02 0.73 3.18 2.70 ;
        RECT  3.02 2.54 3.90 2.70 ;
        RECT  3.62 2.48 3.90 2.76 ;
        RECT  4.76 0.73 5.04 1.01 ;
        RECT  3.98 1.37 4.98 1.53 ;
        RECT  3.98 1.31 4.26 1.59 ;
        RECT  4.82 0.73 4.98 2.18 ;
        RECT  4.76 1.90 5.04 2.18 ;
    END
END DLAHSP8V1_0

MACRO DLAHSP4V1_0
    CLASS CORE ;
    FOREIGN DLAHSP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.99 1.46 2.41 1.74 ;
        END
    END D
    PIN G
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.32 1.40 0.74 1.68 ;
        END
    END G
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 14.88  LAYER ME1  ;
        ANTENNADIFFAREA 7.55  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.95  LAYER ME1  ;
        ANTENNAMAXAREACAR 15.66  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.80 1.84 7.08 2.48 ;
        RECT  6.92 0.60 7.08 2.48 ;
        RECT  6.80 0.60 7.08 1.24 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 14.88  LAYER ME1  ;
        ANTENNADIFFAREA 7.30  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.95  LAYER ME1  ;
        ANTENNAMAXAREACAR 15.66  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.72 1.84 6.04 2.48 ;
        RECT  5.72 0.60 6.04 1.24 ;
        RECT  5.72 0.60 5.88 2.48 ;
        END
    END QB
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 8.00 3.48 ;
        RECT  7.38 2.88 7.82 3.48 ;
        RECT  7.32 1.84 7.60 2.48 ;
        RECT  7.38 1.84 7.54 3.48 ;
        RECT  6.28 1.84 6.56 2.48 ;
        RECT  6.34 1.84 6.50 3.48 ;
        RECT  5.24 1.84 5.52 2.48 ;
        RECT  5.30 1.84 5.46 3.48 ;
        RECT  4.24 1.90 4.52 2.18 ;
        RECT  4.30 1.90 4.46 3.48 ;
        RECT  1.92 1.90 2.20 2.18 ;
        RECT  1.98 1.90 2.14 3.48 ;
        RECT  0.22 1.84 0.50 2.12 ;
        RECT  0.29 1.84 0.45 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 8.00 0.28 ;
        RECT  7.38 -0.28 7.82 0.32 ;
        RECT  7.32 0.60 7.60 1.24 ;
        RECT  7.38 -0.28 7.54 1.24 ;
        RECT  6.28 0.60 6.56 1.24 ;
        RECT  6.34 -0.28 6.50 1.24 ;
        RECT  5.24 0.60 5.52 1.24 ;
        RECT  5.30 -0.28 5.46 1.24 ;
        RECT  4.24 0.73 4.52 1.01 ;
        RECT  4.30 -0.28 4.46 1.01 ;
        RECT  1.92 0.73 2.20 1.01 ;
        RECT  1.98 -0.28 2.14 1.01 ;
        RECT  0.22 0.96 0.50 1.24 ;
        RECT  0.28 -0.28 0.44 1.24 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.74 0.96 1.06 1.24 ;
        RECT  0.90 1.40 1.30 1.68 ;
        RECT  0.90 0.96 1.06 2.12 ;
        RECT  0.74 1.84 1.06 2.12 ;
        RECT  1.40 0.73 1.68 1.01 ;
        RECT  1.46 0.73 1.62 2.18 ;
        RECT  1.34 1.90 1.68 2.18 ;
        RECT  1.34 1.90 1.50 2.76 ;
        RECT  1.22 2.48 1.50 2.76 ;
        RECT  2.44 0.73 2.77 1.01 ;
        RECT  2.61 0.73 2.77 2.18 ;
        RECT  2.44 1.90 2.77 2.18 ;
        RECT  3.48 0.73 3.76 1.01 ;
        RECT  3.54 0.73 3.70 2.18 ;
        RECT  3.48 1.90 3.76 2.18 ;
        RECT  2.96 0.73 3.24 1.01 ;
        RECT  2.96 1.90 3.24 2.18 ;
        RECT  3.02 0.73 3.18 2.70 ;
        RECT  3.02 2.54 3.90 2.70 ;
        RECT  3.62 2.48 3.90 2.76 ;
        RECT  4.76 0.73 5.04 1.01 ;
        RECT  3.98 1.37 4.98 1.53 ;
        RECT  3.98 1.31 4.26 1.59 ;
        RECT  4.82 0.73 4.98 2.18 ;
        RECT  4.76 1.90 5.04 2.18 ;
    END
END DLAHSP4V1_0

MACRO DLAHSP2V1_0
    CLASS CORE ;
    FOREIGN DLAHSP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 12.53  LAYER ME1  ;
        ANTENNADIFFAREA 5.84  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER ME1  ;
        ANTENNAMAXAREACAR 19.78  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.24 1.84 5.52 2.46 ;
        RECT  5.24 0.62 5.52 1.24 ;
        RECT  5.32 0.62 5.48 2.46 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 12.53  LAYER ME1  ;
        ANTENNADIFFAREA 5.84  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER ME1  ;
        ANTENNAMAXAREACAR 19.78  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.28 1.84 6.56 2.46 ;
        RECT  6.28 0.62 6.56 1.24 ;
        RECT  6.34 0.62 6.50 2.46 ;
        RECT  6.12 1.52 6.50 1.68 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.32 1.40 0.74 1.68 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.99 1.46 2.41 1.74 ;
        END
    END D
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 6.80 0.28 ;
        RECT  6.34 -0.28 6.62 0.32 ;
        RECT  5.76 0.62 6.04 1.24 ;
        RECT  5.81 -0.28 5.97 1.24 ;
        RECT  4.24 0.73 4.52 1.01 ;
        RECT  4.30 -0.28 4.46 1.01 ;
        RECT  1.92 0.73 2.20 1.01 ;
        RECT  1.98 -0.28 2.14 1.01 ;
        RECT  0.22 0.96 0.50 1.24 ;
        RECT  0.28 -0.28 0.44 1.24 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 6.80 3.48 ;
        RECT  6.34 2.88 6.62 3.48 ;
        RECT  5.76 1.84 6.04 2.46 ;
        RECT  5.81 1.84 5.97 3.48 ;
        RECT  4.24 1.90 4.52 2.18 ;
        RECT  4.30 1.90 4.46 3.48 ;
        RECT  1.92 1.90 2.20 2.18 ;
        RECT  1.98 1.90 2.14 3.48 ;
        RECT  0.22 1.84 0.50 2.12 ;
        RECT  0.29 1.84 0.45 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.74 0.96 1.06 1.24 ;
        RECT  0.90 1.40 1.30 1.68 ;
        RECT  0.90 0.96 1.06 2.12 ;
        RECT  0.74 1.84 1.06 2.12 ;
        RECT  1.40 0.73 1.68 1.01 ;
        RECT  1.46 0.73 1.62 2.18 ;
        RECT  1.34 1.90 1.68 2.18 ;
        RECT  1.34 1.90 1.50 2.76 ;
        RECT  1.22 2.48 1.50 2.76 ;
        RECT  2.44 0.73 2.77 1.01 ;
        RECT  2.61 0.73 2.77 2.18 ;
        RECT  2.44 1.90 2.77 2.18 ;
        RECT  3.48 0.73 3.76 1.01 ;
        RECT  3.54 0.73 3.70 2.18 ;
        RECT  3.48 1.90 3.76 2.18 ;
        RECT  2.96 0.73 3.24 1.01 ;
        RECT  2.96 1.90 3.24 2.18 ;
        RECT  3.02 0.73 3.18 2.70 ;
        RECT  3.02 2.54 3.90 2.70 ;
        RECT  3.62 2.48 3.90 2.76 ;
        RECT  4.76 0.73 5.04 1.01 ;
        RECT  3.98 1.37 4.98 1.53 ;
        RECT  3.98 1.31 4.26 1.59 ;
        RECT  4.82 0.73 4.98 2.18 ;
        RECT  4.76 1.90 5.04 2.18 ;
    END
END DLAHSP2V1_0

MACRO DLAHSP1V1_0
    CLASS CORE ;
    FOREIGN DLAHSP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.99 1.46 2.41 1.74 ;
        END
    END D
    PIN G
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.32 1.40 0.74 1.68 ;
        END
    END G
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 12.12  LAYER ME1  ;
        ANTENNADIFFAREA 5.11  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.47  LAYER ME1  ;
        ANTENNAMAXAREACAR 25.76  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.28 1.89 6.56 2.17 ;
        RECT  6.28 0.73 6.56 1.01 ;
        RECT  6.34 0.73 6.50 2.17 ;
        RECT  6.12 1.52 6.50 1.68 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 11.82  LAYER ME1  ;
        ANTENNADIFFAREA 5.11  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.47  LAYER ME1  ;
        ANTENNAMAXAREACAR 25.12  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.24 1.89 5.52 2.17 ;
        RECT  5.24 0.73 5.52 1.01 ;
        RECT  5.32 0.73 5.48 2.17 ;
        END
    END QB
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 6.80 3.48 ;
        RECT  6.34 2.88 6.62 3.48 ;
        RECT  5.76 1.89 6.04 2.17 ;
        RECT  5.81 1.89 5.97 3.48 ;
        RECT  4.24 1.90 4.52 2.18 ;
        RECT  4.30 1.90 4.46 3.48 ;
        RECT  1.92 1.90 2.20 2.18 ;
        RECT  1.98 1.90 2.14 3.48 ;
        RECT  0.22 1.84 0.50 2.12 ;
        RECT  0.29 1.84 0.45 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 6.80 0.28 ;
        RECT  6.34 -0.28 6.62 0.32 ;
        RECT  5.76 0.73 6.04 1.01 ;
        RECT  5.81 -0.28 5.97 1.01 ;
        RECT  4.24 0.73 4.52 1.01 ;
        RECT  4.30 -0.28 4.46 1.01 ;
        RECT  1.92 0.73 2.20 1.01 ;
        RECT  1.98 -0.28 2.14 1.01 ;
        RECT  0.22 0.96 0.50 1.24 ;
        RECT  0.28 -0.28 0.44 1.24 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.74 0.96 1.06 1.24 ;
        RECT  0.90 1.40 1.30 1.68 ;
        RECT  0.90 0.96 1.06 2.12 ;
        RECT  0.74 1.84 1.06 2.12 ;
        RECT  1.40 0.73 1.68 1.01 ;
        RECT  1.46 0.73 1.62 2.18 ;
        RECT  1.34 1.90 1.68 2.18 ;
        RECT  1.34 1.90 1.50 2.76 ;
        RECT  1.22 2.48 1.50 2.76 ;
        RECT  2.44 0.73 2.77 1.01 ;
        RECT  2.61 0.73 2.77 2.18 ;
        RECT  2.44 1.90 2.77 2.18 ;
        RECT  3.48 0.73 3.76 1.01 ;
        RECT  3.54 0.73 3.70 2.18 ;
        RECT  3.48 1.90 3.76 2.18 ;
        RECT  2.96 0.73 3.24 1.01 ;
        RECT  2.96 1.90 3.24 2.18 ;
        RECT  3.02 0.73 3.18 2.70 ;
        RECT  3.02 2.54 3.90 2.70 ;
        RECT  3.62 2.48 3.90 2.76 ;
        RECT  4.76 0.73 5.04 1.01 ;
        RECT  3.98 1.37 4.98 1.53 ;
        RECT  3.98 1.31 4.26 1.59 ;
        RECT  4.82 0.73 4.98 2.18 ;
        RECT  4.76 1.90 5.04 2.18 ;
    END
END DLAHSP1V1_0

MACRO DLAHRSP1V1_0
    CLASS CORE ;
    FOREIGN DLAHRSP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 13.90  LAYER ME1  ;
        ANTENNADIFFAREA 5.88  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.47  LAYER ME1  ;
        ANTENNAMAXAREACAR 29.54  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.12 1.89 6.44 2.17 ;
        RECT  6.12 0.73 6.44 1.01 ;
        RECT  6.12 0.73 6.28 2.17 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 13.90  LAYER ME1  ;
        ANTENNADIFFAREA 5.88  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.47  LAYER ME1  ;
        ANTENNAMAXAREACAR 29.54  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.26 1.46 7.50 1.74 ;
        RECT  7.20 1.89 7.48 2.17 ;
        RECT  7.20 0.73 7.48 1.01 ;
        RECT  7.26 0.73 7.42 2.17 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.46 1.40 0.74 1.68 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.86 1.46 3.30 1.74 ;
        END
    END D
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.00 1.46 2.28 1.74 ;
        END
    END RB
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 7.60 0.28 ;
        RECT  7.14 -0.28 7.42 0.32 ;
        RECT  6.68 0.73 6.96 1.01 ;
        RECT  6.73 -0.28 6.89 1.01 ;
        RECT  5.16 0.73 5.44 1.01 ;
        RECT  5.22 -0.28 5.38 1.01 ;
        RECT  2.32 0.70 2.60 0.98 ;
        RECT  2.38 -0.28 2.54 0.98 ;
        RECT  1.84 0.73 2.12 1.01 ;
        RECT  1.90 -0.28 2.06 1.01 ;
        RECT  0.22 0.96 0.50 1.24 ;
        RECT  0.28 -0.28 0.44 1.24 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 7.60 3.48 ;
        RECT  7.14 2.88 7.42 3.48 ;
        RECT  6.68 1.89 6.96 2.17 ;
        RECT  6.73 1.89 6.89 3.48 ;
        RECT  5.16 1.90 5.44 2.18 ;
        RECT  5.22 1.90 5.38 3.48 ;
        RECT  2.84 1.90 3.12 2.18 ;
        RECT  2.90 1.90 3.06 3.48 ;
        RECT  1.84 1.90 2.12 2.18 ;
        RECT  1.90 1.90 2.06 3.48 ;
        RECT  0.22 1.84 0.50 2.12 ;
        RECT  0.29 1.84 0.45 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.74 0.96 1.06 1.24 ;
        RECT  0.90 1.40 1.22 1.68 ;
        RECT  0.90 0.96 1.06 2.12 ;
        RECT  0.74 1.84 1.06 2.12 ;
        RECT  1.32 0.73 1.60 1.01 ;
        RECT  1.38 0.73 1.54 2.18 ;
        RECT  1.26 1.90 1.60 2.18 ;
        RECT  1.26 1.90 1.42 2.76 ;
        RECT  1.14 2.48 1.42 2.76 ;
        RECT  3.40 0.76 3.68 1.04 ;
        RECT  3.53 1.04 3.69 2.18 ;
        RECT  3.36 1.90 3.69 2.18 ;
        RECT  4.46 0.73 4.76 1.01 ;
        RECT  4.46 0.73 4.62 2.18 ;
        RECT  4.40 1.90 4.68 2.18 ;
        RECT  2.76 0.44 4.08 0.60 ;
        RECT  3.92 0.44 4.08 1.04 ;
        RECT  3.92 0.76 4.20 1.04 ;
        RECT  2.76 0.44 2.92 1.30 ;
        RECT  2.44 1.14 2.92 1.30 ;
        RECT  2.44 1.14 2.60 2.18 ;
        RECT  2.32 1.90 2.60 2.18 ;
        RECT  3.88 1.90 4.16 2.18 ;
        RECT  3.94 0.76 4.10 2.70 ;
        RECT  3.94 2.54 4.82 2.70 ;
        RECT  4.54 2.48 4.82 2.76 ;
        RECT  5.68 0.73 5.96 1.01 ;
        RECT  4.90 1.37 5.90 1.53 ;
        RECT  4.90 1.31 5.18 1.59 ;
        RECT  5.74 0.73 5.90 2.18 ;
        RECT  5.68 1.90 5.96 2.18 ;
    END
END DLAHRSP1V1_0

MACRO DFFSZSP8V1_0
    CLASS CORE ;
    FOREIGN DFFSZSP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 21.17  LAYER ME1  ;
        ANTENNADIFFAREA 9.99  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.05  LAYER ME1  ;
        ANTENNAMAXAREACAR 20.23  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.94 1.84 11.22 2.12 ;
        RECT  10.94 0.96 11.22 1.24 ;
        RECT  10.94 0.96 11.10 2.12 ;
        RECT  10.02 1.52 11.10 1.68 ;
        RECT  10.02 1.46 10.34 1.74 ;
        RECT  9.90 1.84 10.18 2.12 ;
        RECT  10.02 0.96 10.18 2.12 ;
        RECT  9.90 0.96 10.18 1.24 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.20  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.85  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.81 1.19 2.25 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  0.91 0.81 1.19 1.09 ;
        END
    END D
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END SEL
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.87  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 12.92  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.06 1.46 2.34 1.74 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.81 2.23 2.25 ;
        RECT  1.95 0.81 2.23 1.09 ;
        END
    END TD
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.21 1.40 3.53 1.80 ;
        END
    END CK
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 12.00 0.28 ;
        RECT  11.52 -0.28 11.82 0.32 ;
        RECT  11.46 0.64 11.74 0.92 ;
        RECT  11.52 -0.28 11.68 0.92 ;
        RECT  10.42 0.64 10.70 0.92 ;
        RECT  10.48 -0.28 10.64 0.92 ;
        RECT  9.38 0.64 9.66 0.92 ;
        RECT  9.44 -0.28 9.60 0.92 ;
        RECT  8.38 0.96 8.66 1.24 ;
        RECT  8.48 -0.28 8.64 1.24 ;
        RECT  5.66 0.72 5.94 1.00 ;
        RECT  5.72 -0.28 5.88 1.00 ;
        RECT  2.95 0.68 3.23 0.96 ;
        RECT  3.01 -0.28 3.17 0.96 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 12.00 3.48 ;
        RECT  11.52 2.88 11.82 3.48 ;
        RECT  11.46 2.16 11.74 2.44 ;
        RECT  11.52 2.16 11.68 3.48 ;
        RECT  10.42 2.16 10.70 2.44 ;
        RECT  10.48 2.16 10.64 3.48 ;
        RECT  9.38 2.16 9.66 2.44 ;
        RECT  9.44 2.16 9.60 3.48 ;
        RECT  8.38 2.62 8.66 3.48 ;
        RECT  5.81 1.92 6.09 2.20 ;
        RECT  5.87 1.92 6.03 3.48 ;
        RECT  2.71 2.62 2.99 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  1.55 1.97 1.71 2.58 ;
        RECT  1.55 2.42 2.37 2.58 ;
        RECT  2.09 2.41 2.37 2.69 ;
        RECT  3.47 0.68 3.85 0.96 ;
        RECT  3.69 1.22 3.97 1.50 ;
        RECT  3.69 0.68 3.85 2.25 ;
        RECT  3.47 1.97 3.85 2.25 ;
        RECT  2.43 0.68 2.71 0.96 ;
        RECT  4.01 0.72 4.29 1.00 ;
        RECT  2.55 0.68 2.71 2.25 ;
        RECT  2.43 1.97 2.71 2.25 ;
        RECT  4.13 0.72 4.29 2.20 ;
        RECT  2.43 2.09 3.31 2.25 ;
        RECT  3.15 2.09 3.31 2.57 ;
        RECT  4.01 1.92 4.17 2.57 ;
        RECT  3.15 2.41 4.17 2.57 ;
        RECT  5.09 0.72 5.39 1.00 ;
        RECT  5.09 0.72 5.25 2.20 ;
        RECT  5.05 1.92 5.33 2.20 ;
        RECT  4.53 0.72 4.81 1.00 ;
        RECT  5.89 1.48 6.17 1.76 ;
        RECT  5.49 1.60 6.17 1.76 ;
        RECT  4.59 0.72 4.75 2.20 ;
        RECT  4.53 1.92 4.81 2.20 ;
        RECT  4.65 1.92 4.81 2.52 ;
        RECT  5.49 1.60 5.65 2.52 ;
        RECT  4.65 2.36 5.65 2.52 ;
        RECT  6.18 0.72 6.49 1.00 ;
        RECT  5.41 1.16 6.49 1.32 ;
        RECT  5.41 1.16 5.69 1.44 ;
        RECT  6.33 0.72 6.49 2.20 ;
        RECT  6.33 1.92 6.61 2.20 ;
        RECT  6.86 0.44 8.32 0.60 ;
        RECT  8.04 0.44 8.32 0.80 ;
        RECT  6.74 0.76 7.02 1.04 ;
        RECT  6.86 0.44 7.02 2.20 ;
        RECT  6.85 1.92 7.13 2.20 ;
        RECT  7.86 0.96 8.14 1.24 ;
        RECT  7.86 1.46 8.86 1.62 ;
        RECT  8.58 1.40 8.86 1.68 ;
        RECT  7.86 0.96 8.02 2.12 ;
        RECT  7.86 1.84 8.14 2.12 ;
        RECT  7.26 0.76 7.54 1.04 ;
        RECT  8.90 0.96 9.18 1.24 ;
        RECT  8.90 1.84 9.18 2.12 ;
        RECT  7.38 0.76 7.54 2.20 ;
        RECT  7.37 1.92 7.65 2.20 ;
        RECT  7.49 1.92 7.65 2.44 ;
        RECT  9.02 0.96 9.18 2.44 ;
        RECT  7.49 2.28 9.18 2.44 ;
    END
END DFFSZSP8V1_0

MACRO DFFSZSP4V1_0
    CLASS CORE ;
    FOREIGN DFFSZSP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 18.89  LAYER ME1  ;
        ANTENNADIFFAREA 8.44  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.76  LAYER ME1  ;
        ANTENNAMAXAREACAR 24.90  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.02 1.46 10.34 1.74 ;
        RECT  9.90 1.84 10.18 2.12 ;
        RECT  10.02 0.96 10.18 2.12 ;
        RECT  9.90 0.96 10.18 1.24 ;
        END
    END Q
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.21 1.40 3.53 1.80 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.87  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 12.92  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.06 1.46 2.34 1.74 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.81 2.23 2.25 ;
        RECT  1.95 0.81 2.23 1.09 ;
        END
    END TD
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END SEL
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.20  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.85  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.81 1.19 2.25 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  0.91 0.81 1.19 1.09 ;
        END
    END D
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 10.80 0.28 ;
        RECT  10.42 0.64 10.70 0.92 ;
        RECT  10.48 -0.28 10.64 0.92 ;
        RECT  10.34 -0.28 10.64 0.32 ;
        RECT  9.38 0.64 9.66 0.92 ;
        RECT  9.44 -0.28 9.60 0.92 ;
        RECT  8.38 0.96 8.66 1.24 ;
        RECT  8.48 -0.28 8.64 1.24 ;
        RECT  5.66 0.72 5.94 1.00 ;
        RECT  5.72 -0.28 5.88 1.00 ;
        RECT  2.95 0.68 3.23 0.96 ;
        RECT  3.01 -0.28 3.17 0.96 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 10.80 3.48 ;
        RECT  10.42 2.16 10.70 2.44 ;
        RECT  10.34 2.88 10.64 3.48 ;
        RECT  10.48 2.16 10.64 3.48 ;
        RECT  9.38 2.16 9.66 2.44 ;
        RECT  9.44 2.16 9.60 3.48 ;
        RECT  8.38 2.62 8.66 3.48 ;
        RECT  5.81 1.92 6.09 2.20 ;
        RECT  5.87 1.92 6.03 3.48 ;
        RECT  2.71 2.62 2.99 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  1.55 1.97 1.71 2.58 ;
        RECT  1.55 2.42 2.37 2.58 ;
        RECT  2.09 2.41 2.37 2.69 ;
        RECT  3.47 0.68 3.85 0.96 ;
        RECT  3.69 1.22 3.97 1.50 ;
        RECT  3.69 0.68 3.85 2.25 ;
        RECT  3.47 1.97 3.85 2.25 ;
        RECT  2.43 0.68 2.71 0.96 ;
        RECT  4.01 0.72 4.29 1.00 ;
        RECT  2.55 0.68 2.71 2.25 ;
        RECT  2.43 1.97 2.71 2.25 ;
        RECT  4.13 0.72 4.29 2.20 ;
        RECT  2.43 2.09 3.31 2.25 ;
        RECT  3.15 2.09 3.31 2.57 ;
        RECT  4.01 1.92 4.17 2.57 ;
        RECT  3.15 2.41 4.17 2.57 ;
        RECT  5.09 0.72 5.39 1.00 ;
        RECT  5.09 0.72 5.25 2.20 ;
        RECT  5.05 1.92 5.33 2.20 ;
        RECT  4.53 0.72 4.81 1.00 ;
        RECT  5.89 1.48 6.17 1.76 ;
        RECT  5.49 1.60 6.17 1.76 ;
        RECT  4.59 0.72 4.75 2.20 ;
        RECT  4.53 1.92 4.81 2.20 ;
        RECT  4.65 1.92 4.81 2.52 ;
        RECT  5.49 1.60 5.65 2.52 ;
        RECT  4.65 2.36 5.65 2.52 ;
        RECT  6.18 0.72 6.49 1.00 ;
        RECT  5.41 1.16 6.49 1.32 ;
        RECT  5.41 1.16 5.69 1.44 ;
        RECT  6.33 0.72 6.49 2.20 ;
        RECT  6.33 1.92 6.61 2.20 ;
        RECT  6.86 0.44 8.32 0.60 ;
        RECT  8.04 0.44 8.32 0.80 ;
        RECT  6.74 0.76 7.02 1.04 ;
        RECT  6.86 0.44 7.02 2.20 ;
        RECT  6.85 1.92 7.13 2.20 ;
        RECT  7.86 0.96 8.14 1.24 ;
        RECT  7.86 1.46 8.86 1.62 ;
        RECT  8.58 1.40 8.86 1.68 ;
        RECT  7.86 0.96 8.02 2.12 ;
        RECT  7.86 1.84 8.14 2.12 ;
        RECT  7.26 0.76 7.54 1.04 ;
        RECT  8.90 0.96 9.18 1.24 ;
        RECT  8.90 1.84 9.18 2.12 ;
        RECT  7.38 0.76 7.54 2.20 ;
        RECT  7.37 1.92 7.65 2.20 ;
        RECT  7.49 1.92 7.65 2.44 ;
        RECT  9.02 0.96 9.18 2.44 ;
        RECT  7.49 2.28 9.18 2.44 ;
    END
END DFFSZSP4V1_0

MACRO DFFSZSP2V1_0
    CLASS CORE ;
    FOREIGN DFFSZSP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.20  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.85  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.81 1.19 2.25 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  0.91 0.81 1.19 1.09 ;
        END
    END D
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END SEL
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.87  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 12.92  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.06 1.46 2.34 1.74 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.81 2.23 2.25 ;
        RECT  1.95 0.81 2.23 1.09 ;
        END
    END TD
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.21 1.40 3.53 1.80 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 18.16  LAYER ME1  ;
        ANTENNADIFFAREA 7.84  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.61  LAYER ME1  ;
        ANTENNAMAXAREACAR 29.56  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.05 1.46 10.32 1.74 ;
        RECT  9.93 1.84 10.21 2.12 ;
        RECT  10.05 0.96 10.21 2.12 ;
        RECT  9.93 0.96 10.21 1.24 ;
        END
    END Q
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 10.40 3.48 ;
        RECT  9.94 2.88 10.22 3.48 ;
        RECT  9.41 2.16 9.69 2.44 ;
        RECT  9.47 2.16 9.63 3.48 ;
        RECT  8.41 2.62 8.69 3.48 ;
        RECT  5.81 1.92 6.09 2.20 ;
        RECT  5.87 1.92 6.03 3.48 ;
        RECT  2.71 2.62 2.99 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 10.40 0.28 ;
        RECT  9.94 -0.28 10.22 0.32 ;
        RECT  9.41 0.64 9.69 0.92 ;
        RECT  9.47 -0.28 9.63 0.92 ;
        RECT  8.41 0.96 8.69 1.24 ;
        RECT  8.51 -0.28 8.67 1.24 ;
        RECT  5.69 0.72 5.97 1.00 ;
        RECT  5.75 -0.28 5.91 1.00 ;
        RECT  2.95 0.68 3.23 0.96 ;
        RECT  3.01 -0.28 3.17 0.96 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  1.55 1.97 1.71 2.58 ;
        RECT  1.55 2.42 2.37 2.58 ;
        RECT  2.09 2.41 2.37 2.69 ;
        RECT  3.47 0.68 3.85 0.96 ;
        RECT  3.69 1.22 3.97 1.50 ;
        RECT  3.69 0.68 3.85 2.25 ;
        RECT  3.47 1.97 3.85 2.25 ;
        RECT  2.43 0.68 2.71 0.96 ;
        RECT  4.01 0.72 4.29 1.00 ;
        RECT  2.55 0.68 2.71 2.25 ;
        RECT  2.43 1.97 2.71 2.25 ;
        RECT  4.13 0.72 4.29 2.20 ;
        RECT  2.43 2.09 3.31 2.25 ;
        RECT  3.15 2.09 3.31 2.57 ;
        RECT  4.01 1.92 4.17 2.57 ;
        RECT  3.15 2.41 4.17 2.57 ;
        RECT  5.09 0.72 5.40 1.00 ;
        RECT  5.09 0.72 5.25 2.20 ;
        RECT  5.05 1.92 5.33 2.20 ;
        RECT  4.53 0.72 4.81 1.00 ;
        RECT  5.89 1.48 6.17 1.76 ;
        RECT  5.49 1.60 6.17 1.76 ;
        RECT  4.59 0.72 4.75 2.20 ;
        RECT  4.53 1.92 4.81 2.20 ;
        RECT  4.65 1.92 4.81 2.52 ;
        RECT  5.49 1.60 5.65 2.52 ;
        RECT  4.65 2.36 5.65 2.52 ;
        RECT  6.21 0.72 6.49 1.00 ;
        RECT  5.41 1.16 6.49 1.32 ;
        RECT  5.41 1.16 5.69 1.44 ;
        RECT  6.33 0.72 6.49 2.20 ;
        RECT  6.33 1.92 6.61 2.20 ;
        RECT  6.89 0.44 8.35 0.60 ;
        RECT  8.07 0.44 8.35 0.80 ;
        RECT  6.77 0.76 7.05 1.04 ;
        RECT  6.89 0.44 7.05 2.20 ;
        RECT  6.85 1.92 7.13 2.20 ;
        RECT  7.89 0.96 8.17 1.24 ;
        RECT  7.89 1.46 8.89 1.62 ;
        RECT  8.61 1.40 8.89 1.68 ;
        RECT  7.89 0.96 8.05 2.12 ;
        RECT  7.89 1.84 8.17 2.12 ;
        RECT  7.29 0.76 7.57 1.04 ;
        RECT  8.93 0.96 9.21 1.24 ;
        RECT  8.93 1.84 9.21 2.12 ;
        RECT  7.41 0.76 7.57 2.20 ;
        RECT  7.37 1.92 7.65 2.20 ;
        RECT  7.49 1.92 7.65 2.44 ;
        RECT  9.05 0.96 9.21 2.44 ;
        RECT  7.49 2.28 9.21 2.44 ;
    END
END DFFSZSP2V1_0

MACRO DFFSZSP1V1_0
    CLASS CORE ;
    FOREIGN DFFSZSP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 18.26  LAYER ME1  ;
        ANTENNADIFFAREA 7.40  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.54  LAYER ME1  ;
        ANTENNAMAXAREACAR 33.97  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.05 1.46 10.32 1.74 ;
        RECT  9.93 1.84 10.21 2.12 ;
        RECT  10.05 0.96 10.21 2.12 ;
        RECT  9.93 0.96 10.21 1.24 ;
        END
    END Q
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.21 1.40 3.53 1.80 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.20  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.85  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.81 1.19 2.25 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  0.91 0.81 1.19 1.09 ;
        END
    END D
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.87  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 12.92  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.06 1.46 2.34 1.74 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.81 2.23 2.25 ;
        RECT  1.95 0.81 2.23 1.09 ;
        END
    END TD
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END SEL
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 10.40 0.28 ;
        RECT  9.94 -0.28 10.22 0.32 ;
        RECT  9.41 0.96 9.69 1.24 ;
        RECT  9.47 -0.28 9.63 1.24 ;
        RECT  8.41 0.96 8.69 1.24 ;
        RECT  8.51 -0.28 8.67 1.24 ;
        RECT  5.69 0.72 5.97 1.00 ;
        RECT  5.75 -0.28 5.91 1.00 ;
        RECT  2.95 0.68 3.23 0.96 ;
        RECT  3.01 -0.28 3.17 0.96 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 10.40 3.48 ;
        RECT  9.94 2.88 10.22 3.48 ;
        RECT  9.41 1.84 9.69 2.12 ;
        RECT  9.47 1.84 9.63 3.48 ;
        RECT  8.41 2.62 8.69 3.48 ;
        RECT  5.81 1.92 6.09 2.20 ;
        RECT  5.87 1.92 6.03 3.48 ;
        RECT  2.71 2.62 2.99 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  1.55 1.97 1.71 2.58 ;
        RECT  1.55 2.42 2.37 2.58 ;
        RECT  2.09 2.41 2.37 2.69 ;
        RECT  3.47 0.68 3.85 0.96 ;
        RECT  3.69 1.22 3.97 1.50 ;
        RECT  3.69 0.68 3.85 2.25 ;
        RECT  3.47 1.97 3.85 2.25 ;
        RECT  2.43 0.68 2.71 0.96 ;
        RECT  4.01 0.72 4.29 1.00 ;
        RECT  2.55 0.68 2.71 2.25 ;
        RECT  2.43 1.97 2.71 2.25 ;
        RECT  4.13 0.72 4.29 2.20 ;
        RECT  2.43 2.09 3.31 2.25 ;
        RECT  3.15 2.09 3.31 2.57 ;
        RECT  4.01 1.92 4.17 2.57 ;
        RECT  3.15 2.41 4.17 2.57 ;
        RECT  5.09 0.72 5.40 1.00 ;
        RECT  5.09 0.72 5.25 2.20 ;
        RECT  5.05 1.92 5.33 2.20 ;
        RECT  4.53 0.72 4.81 1.00 ;
        RECT  5.89 1.48 6.17 1.76 ;
        RECT  5.49 1.60 6.17 1.76 ;
        RECT  4.59 0.72 4.75 2.20 ;
        RECT  4.53 1.92 4.81 2.20 ;
        RECT  4.65 1.92 4.81 2.52 ;
        RECT  5.49 1.60 5.65 2.52 ;
        RECT  4.65 2.36 5.65 2.52 ;
        RECT  6.21 0.72 6.49 1.00 ;
        RECT  5.41 1.16 6.49 1.32 ;
        RECT  5.41 1.16 5.69 1.44 ;
        RECT  6.33 0.72 6.49 2.20 ;
        RECT  6.33 1.92 6.61 2.20 ;
        RECT  6.89 0.44 8.35 0.60 ;
        RECT  8.07 0.44 8.35 0.80 ;
        RECT  6.77 0.76 7.05 1.04 ;
        RECT  6.89 0.44 7.05 2.20 ;
        RECT  6.85 1.92 7.13 2.20 ;
        RECT  7.89 0.96 8.17 1.24 ;
        RECT  7.89 1.46 8.89 1.62 ;
        RECT  8.61 1.40 8.89 1.68 ;
        RECT  7.89 0.96 8.05 2.12 ;
        RECT  7.89 1.84 8.17 2.12 ;
        RECT  7.29 0.76 7.57 1.04 ;
        RECT  8.93 0.96 9.21 1.24 ;
        RECT  8.93 1.84 9.21 2.12 ;
        RECT  7.41 0.76 7.57 2.20 ;
        RECT  7.37 1.92 7.65 2.20 ;
        RECT  7.49 1.92 7.65 2.44 ;
        RECT  9.05 0.96 9.21 2.44 ;
        RECT  7.49 2.28 9.21 2.44 ;
    END
END DFFSZSP1V1_0

MACRO DFFSSZSP8V1_0
    CLASS CORE ;
    FOREIGN DFFSSZSP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 26.96  LAYER ME1  ;
        ANTENNADIFFAREA 12.39  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.05  LAYER ME1  ;
        ANTENNAMAXAREACAR 25.77  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.17 1.90 13.45 2.50 ;
        RECT  13.17 0.64 13.45 1.24 ;
        RECT  13.17 0.64 13.33 2.50 ;
        RECT  12.06 1.52 13.33 1.68 ;
        RECT  12.13 1.90 12.41 2.50 ;
        RECT  12.13 0.64 12.41 1.24 ;
        RECT  12.13 0.64 12.34 2.50 ;
        RECT  12.06 1.46 12.34 1.74 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.52 1.40 9.94 1.68 ;
        END
    END SB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.24 1.40 3.54 1.76 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.87  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 12.90  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.06 1.46 2.34 1.74 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.81 2.23 2.25 ;
        RECT  1.95 0.81 2.23 1.09 ;
        END
    END TD
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END SEL
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.20  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.83  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.81 1.19 2.25 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  0.91 0.81 1.19 1.09 ;
        END
    END D
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 14.40 0.28 ;
        RECT  13.78 -0.28 14.22 0.32 ;
        RECT  13.69 0.64 13.97 1.24 ;
        RECT  13.78 -0.28 13.94 1.24 ;
        RECT  12.65 0.64 12.93 1.24 ;
        RECT  12.71 -0.28 12.87 1.24 ;
        RECT  11.61 0.64 11.89 1.24 ;
        RECT  11.67 -0.28 11.83 1.24 ;
        RECT  10.61 0.88 10.89 1.16 ;
        RECT  10.67 -0.28 10.83 1.16 ;
        RECT  9.13 -0.28 9.41 0.68 ;
        RECT  2.71 -0.28 2.99 0.68 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 14.40 3.48 ;
        RECT  13.78 2.88 14.22 3.48 ;
        RECT  13.69 1.90 13.97 2.50 ;
        RECT  13.78 1.90 13.94 3.48 ;
        RECT  12.65 1.90 12.93 2.50 ;
        RECT  12.71 1.90 12.87 3.48 ;
        RECT  11.61 1.90 11.89 2.50 ;
        RECT  11.67 1.90 11.83 3.48 ;
        RECT  10.37 2.40 10.65 3.48 ;
        RECT  9.57 1.84 9.85 2.12 ;
        RECT  9.63 1.84 9.79 3.48 ;
        RECT  8.57 1.84 8.85 2.12 ;
        RECT  8.63 1.84 8.79 3.48 ;
        RECT  7.57 1.84 7.85 2.12 ;
        RECT  7.67 1.84 7.83 3.48 ;
        RECT  2.71 2.52 2.99 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  1.55 1.97 1.71 2.57 ;
        RECT  1.55 2.41 2.37 2.57 ;
        RECT  2.09 2.41 2.37 2.69 ;
        RECT  3.47 0.96 3.86 1.24 ;
        RECT  3.70 1.46 4.02 1.74 ;
        RECT  3.70 0.96 3.86 2.20 ;
        RECT  3.47 1.92 3.86 2.20 ;
        RECT  4.07 0.44 4.35 0.72 ;
        RECT  3.15 0.56 4.35 0.72 ;
        RECT  3.15 0.56 3.31 1.12 ;
        RECT  2.43 0.96 3.31 1.12 ;
        RECT  2.43 0.96 2.71 1.24 ;
        RECT  2.55 0.96 2.71 2.20 ;
        RECT  2.43 1.92 2.71 2.20 ;
        RECT  2.43 2.04 3.31 2.20 ;
        RECT  3.15 2.04 3.31 2.64 ;
        RECT  3.15 2.48 4.25 2.64 ;
        RECT  3.97 2.48 4.25 2.76 ;
        RECT  5.59 0.76 5.91 1.04 ;
        RECT  5.59 0.76 5.75 2.00 ;
        RECT  5.25 1.84 6.29 2.00 ;
        RECT  5.25 1.84 5.53 2.12 ;
        RECT  6.01 1.84 6.29 2.12 ;
        RECT  6.15 0.76 6.43 1.04 ;
        RECT  6.27 0.76 6.43 1.36 ;
        RECT  7.11 1.08 7.39 1.36 ;
        RECT  6.27 1.20 7.39 1.36 ;
        RECT  6.53 1.20 6.69 2.12 ;
        RECT  6.53 1.84 6.81 2.12 ;
        RECT  4.63 0.86 4.91 1.14 ;
        RECT  4.07 0.98 4.91 1.14 ;
        RECT  4.07 0.96 4.35 1.24 ;
        RECT  4.29 0.98 4.45 2.12 ;
        RECT  4.41 1.84 4.57 2.44 ;
        RECT  4.41 2.28 7.51 2.44 ;
        RECT  7.23 2.28 7.51 2.56 ;
        RECT  6.67 0.76 7.95 0.92 ;
        RECT  6.67 0.76 6.95 1.04 ;
        RECT  7.67 0.76 7.95 1.16 ;
        RECT  7.67 0.76 7.83 1.68 ;
        RECT  8.71 1.40 8.99 1.68 ;
        RECT  7.25 1.52 8.99 1.68 ;
        RECT  8.01 1.52 8.17 2.12 ;
        RECT  7.25 1.52 7.41 2.12 ;
        RECT  7.05 1.84 7.41 2.12 ;
        RECT  8.01 1.84 8.37 2.12 ;
        RECT  5.27 0.44 8.87 0.60 ;
        RECT  8.71 0.44 8.87 1.04 ;
        RECT  8.71 0.88 9.37 1.04 ;
        RECT  5.27 0.44 5.43 1.14 ;
        RECT  9.09 0.88 9.37 1.16 ;
        RECT  5.15 0.86 5.31 1.46 ;
        RECT  4.93 1.30 5.31 1.46 ;
        RECT  9.15 0.88 9.31 2.12 ;
        RECT  4.93 1.30 5.09 2.12 ;
        RECT  4.81 1.84 5.09 2.12 ;
        RECT  9.09 1.84 9.37 2.12 ;
        RECT  9.71 0.88 9.99 1.16 ;
        RECT  9.71 1.00 10.26 1.16 ;
        RECT  10.10 1.00 10.26 2.12 ;
        RECT  10.09 1.84 10.37 2.12 ;
        RECT  10.09 1.96 10.97 2.12 ;
        RECT  10.81 1.96 10.97 2.64 ;
        RECT  10.81 2.48 11.44 2.64 ;
        RECT  11.16 2.48 11.44 2.76 ;
        RECT  11.13 0.88 11.41 1.16 ;
        RECT  10.43 1.46 11.55 1.62 ;
        RECT  10.43 1.40 10.71 1.68 ;
        RECT  11.25 1.40 11.55 1.68 ;
        RECT  11.25 0.88 11.41 2.12 ;
        RECT  11.13 1.84 11.41 2.12 ;
    END
END DFFSSZSP8V1_0

MACRO DFFSSZSP4V1_0
    CLASS CORE ;
    FOREIGN DFFSSZSP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 13.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.20  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.83  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.81 1.19 2.25 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  0.91 0.81 1.19 1.09 ;
        END
    END D
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END SEL
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.87  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 12.90  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.06 1.46 2.34 1.74 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.81 2.23 2.25 ;
        RECT  1.95 0.81 2.23 1.09 ;
        END
    END TD
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.24 1.40 3.54 1.76 ;
        END
    END CK
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.52 1.40 9.94 1.68 ;
        END
    END SB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 24.57  LAYER ME1  ;
        ANTENNADIFFAREA 10.57  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.76  LAYER ME1  ;
        ANTENNAMAXAREACAR 32.40  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.13 1.90 12.41 2.50 ;
        RECT  12.13 0.64 12.41 1.24 ;
        RECT  12.13 0.64 12.34 2.50 ;
        RECT  12.06 1.46 12.34 1.74 ;
        END
    END Q
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 13.20 3.48 ;
        RECT  12.71 2.88 13.02 3.48 ;
        RECT  12.65 1.90 12.93 2.50 ;
        RECT  12.71 1.90 12.87 3.48 ;
        RECT  11.61 1.90 11.89 2.50 ;
        RECT  11.67 1.90 11.83 3.48 ;
        RECT  10.37 2.40 10.65 3.48 ;
        RECT  9.57 1.84 9.85 2.12 ;
        RECT  9.63 1.84 9.79 3.48 ;
        RECT  8.57 1.84 8.85 2.12 ;
        RECT  8.63 1.84 8.79 3.48 ;
        RECT  7.57 1.84 7.85 2.12 ;
        RECT  7.67 1.84 7.83 3.48 ;
        RECT  2.71 2.52 2.99 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 13.20 0.28 ;
        RECT  12.71 -0.28 13.02 0.32 ;
        RECT  12.65 0.64 12.93 1.24 ;
        RECT  12.71 -0.28 12.87 1.24 ;
        RECT  11.61 0.64 11.89 1.24 ;
        RECT  11.67 -0.28 11.83 1.24 ;
        RECT  10.61 0.88 10.89 1.16 ;
        RECT  10.67 -0.28 10.83 1.16 ;
        RECT  9.13 -0.28 9.41 0.68 ;
        RECT  2.71 -0.28 2.99 0.68 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  1.55 1.97 1.71 2.57 ;
        RECT  1.55 2.41 2.37 2.57 ;
        RECT  2.09 2.41 2.37 2.69 ;
        RECT  3.47 0.96 3.86 1.24 ;
        RECT  3.70 1.46 4.02 1.74 ;
        RECT  3.70 0.96 3.86 2.20 ;
        RECT  3.47 1.92 3.86 2.20 ;
        RECT  4.07 0.44 4.35 0.72 ;
        RECT  3.15 0.56 4.35 0.72 ;
        RECT  3.15 0.56 3.31 1.12 ;
        RECT  2.43 0.96 3.31 1.12 ;
        RECT  2.43 0.96 2.71 1.24 ;
        RECT  2.55 0.96 2.71 2.20 ;
        RECT  2.43 1.92 2.71 2.20 ;
        RECT  2.43 2.04 3.31 2.20 ;
        RECT  3.15 2.04 3.31 2.64 ;
        RECT  3.15 2.48 4.25 2.64 ;
        RECT  3.97 2.48 4.25 2.76 ;
        RECT  5.59 0.76 5.91 1.04 ;
        RECT  5.59 0.76 5.75 2.00 ;
        RECT  5.25 1.84 6.29 2.00 ;
        RECT  5.25 1.84 5.53 2.12 ;
        RECT  6.01 1.84 6.29 2.12 ;
        RECT  6.15 0.76 6.43 1.04 ;
        RECT  6.27 0.76 6.43 1.36 ;
        RECT  7.11 1.08 7.39 1.36 ;
        RECT  6.27 1.20 7.39 1.36 ;
        RECT  6.53 1.20 6.69 2.12 ;
        RECT  6.53 1.84 6.81 2.12 ;
        RECT  4.63 0.86 4.91 1.14 ;
        RECT  4.07 0.98 4.91 1.14 ;
        RECT  4.07 0.96 4.35 1.24 ;
        RECT  4.29 0.98 4.45 2.12 ;
        RECT  4.41 1.84 4.57 2.44 ;
        RECT  4.41 2.28 7.51 2.44 ;
        RECT  7.23 2.28 7.51 2.56 ;
        RECT  6.67 0.76 7.95 0.92 ;
        RECT  6.67 0.76 6.95 1.04 ;
        RECT  7.67 0.76 7.95 1.16 ;
        RECT  7.67 0.76 7.83 1.68 ;
        RECT  8.71 1.40 8.99 1.68 ;
        RECT  7.25 1.52 8.99 1.68 ;
        RECT  8.01 1.52 8.17 2.12 ;
        RECT  7.25 1.52 7.41 2.12 ;
        RECT  7.05 1.84 7.41 2.12 ;
        RECT  8.01 1.84 8.37 2.12 ;
        RECT  5.27 0.44 8.87 0.60 ;
        RECT  8.71 0.44 8.87 1.04 ;
        RECT  8.71 0.88 9.37 1.04 ;
        RECT  5.27 0.44 5.43 1.14 ;
        RECT  9.09 0.88 9.37 1.16 ;
        RECT  5.15 0.86 5.31 1.46 ;
        RECT  4.93 1.30 5.31 1.46 ;
        RECT  9.15 0.88 9.31 2.12 ;
        RECT  4.93 1.30 5.09 2.12 ;
        RECT  4.81 1.84 5.09 2.12 ;
        RECT  9.09 1.84 9.37 2.12 ;
        RECT  9.71 0.88 9.99 1.16 ;
        RECT  9.71 1.00 10.26 1.16 ;
        RECT  10.10 1.00 10.26 2.12 ;
        RECT  10.09 1.84 10.37 2.12 ;
        RECT  10.09 1.96 10.97 2.12 ;
        RECT  10.81 1.96 10.97 2.64 ;
        RECT  10.81 2.48 11.44 2.64 ;
        RECT  11.16 2.48 11.44 2.76 ;
        RECT  11.13 0.88 11.41 1.16 ;
        RECT  10.43 1.46 11.55 1.62 ;
        RECT  10.43 1.40 10.71 1.68 ;
        RECT  11.25 1.40 11.55 1.68 ;
        RECT  11.25 0.88 11.41 2.12 ;
        RECT  11.13 1.84 11.41 2.12 ;
    END
END DFFSSZSP4V1_0

MACRO DFFSSZSP2V1_0
    CLASS CORE ;
    FOREIGN DFFSSZSP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 23.75  LAYER ME1  ;
        ANTENNADIFFAREA 9.96  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.61  LAYER ME1  ;
        ANTENNAMAXAREACAR 38.65  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.73 1.46 12.34 1.74 ;
        RECT  11.61 1.90 11.89 2.50 ;
        RECT  11.73 0.64 11.89 2.50 ;
        RECT  11.61 0.64 11.89 1.24 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.52 1.40 9.94 1.68 ;
        END
    END SB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.24 1.40 3.54 1.76 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.87  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 12.90  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.06 1.46 2.34 1.74 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.81 2.23 2.25 ;
        RECT  1.95 0.81 2.23 1.09 ;
        END
    END TD
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END SEL
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.20  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.83  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.81 1.19 2.25 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  0.91 0.81 1.19 1.09 ;
        END
    END D
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 12.80 0.28 ;
        RECT  12.19 -0.28 12.62 0.32 ;
        RECT  12.13 0.64 12.41 1.24 ;
        RECT  12.19 -0.28 12.35 1.24 ;
        RECT  10.61 0.88 10.89 1.16 ;
        RECT  10.67 -0.28 10.83 1.16 ;
        RECT  9.13 -0.28 9.41 0.68 ;
        RECT  2.71 -0.28 2.99 0.68 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 12.80 3.48 ;
        RECT  12.19 2.88 12.62 3.48 ;
        RECT  12.13 1.90 12.41 2.50 ;
        RECT  12.19 1.90 12.35 3.48 ;
        RECT  10.37 2.40 10.65 3.48 ;
        RECT  9.57 1.84 9.85 2.12 ;
        RECT  9.63 1.84 9.79 3.48 ;
        RECT  8.57 1.84 8.85 2.12 ;
        RECT  8.63 1.84 8.79 3.48 ;
        RECT  7.57 1.84 7.85 2.12 ;
        RECT  7.67 1.84 7.83 3.48 ;
        RECT  2.71 2.52 2.99 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  1.55 1.97 1.71 2.57 ;
        RECT  1.55 2.41 2.37 2.57 ;
        RECT  2.09 2.41 2.37 2.69 ;
        RECT  3.47 0.96 3.86 1.24 ;
        RECT  3.70 1.46 4.02 1.74 ;
        RECT  3.70 0.96 3.86 2.20 ;
        RECT  3.47 1.92 3.86 2.20 ;
        RECT  4.07 0.44 4.35 0.72 ;
        RECT  3.15 0.56 4.35 0.72 ;
        RECT  3.15 0.56 3.31 1.12 ;
        RECT  2.43 0.96 3.31 1.12 ;
        RECT  2.43 0.96 2.71 1.24 ;
        RECT  2.55 0.96 2.71 2.20 ;
        RECT  2.43 1.92 2.71 2.20 ;
        RECT  2.43 2.04 3.31 2.20 ;
        RECT  3.15 2.04 3.31 2.64 ;
        RECT  3.15 2.48 4.25 2.64 ;
        RECT  3.97 2.48 4.25 2.76 ;
        RECT  5.59 0.76 5.91 1.04 ;
        RECT  5.59 0.76 5.75 2.00 ;
        RECT  5.25 1.84 6.29 2.00 ;
        RECT  5.25 1.84 5.53 2.12 ;
        RECT  6.01 1.84 6.29 2.12 ;
        RECT  6.15 0.76 6.43 1.04 ;
        RECT  6.27 0.76 6.43 1.36 ;
        RECT  7.11 1.08 7.39 1.36 ;
        RECT  6.27 1.20 7.39 1.36 ;
        RECT  6.53 1.20 6.69 2.12 ;
        RECT  6.53 1.84 6.81 2.12 ;
        RECT  4.63 0.86 4.91 1.14 ;
        RECT  4.07 0.98 4.91 1.14 ;
        RECT  4.07 0.96 4.35 1.24 ;
        RECT  4.29 0.98 4.45 2.12 ;
        RECT  4.41 1.84 4.57 2.44 ;
        RECT  4.41 2.28 7.51 2.44 ;
        RECT  7.23 2.28 7.51 2.56 ;
        RECT  6.67 0.76 7.95 0.92 ;
        RECT  6.67 0.76 6.95 1.04 ;
        RECT  7.67 0.76 7.95 1.16 ;
        RECT  7.67 0.76 7.83 1.68 ;
        RECT  8.71 1.40 8.99 1.68 ;
        RECT  7.25 1.52 8.99 1.68 ;
        RECT  8.01 1.52 8.17 2.12 ;
        RECT  7.25 1.52 7.41 2.12 ;
        RECT  7.05 1.84 7.41 2.12 ;
        RECT  8.01 1.84 8.37 2.12 ;
        RECT  5.27 0.44 8.87 0.60 ;
        RECT  8.71 0.44 8.87 1.04 ;
        RECT  8.71 0.88 9.37 1.04 ;
        RECT  5.27 0.44 5.43 1.14 ;
        RECT  9.09 0.88 9.37 1.16 ;
        RECT  5.15 0.86 5.31 1.46 ;
        RECT  4.93 1.30 5.31 1.46 ;
        RECT  9.15 0.88 9.31 2.12 ;
        RECT  4.93 1.30 5.09 2.12 ;
        RECT  4.81 1.84 5.09 2.12 ;
        RECT  9.09 1.84 9.37 2.12 ;
        RECT  9.71 0.88 9.99 1.16 ;
        RECT  9.71 1.00 10.26 1.16 ;
        RECT  10.10 1.00 10.26 2.12 ;
        RECT  10.09 1.84 10.37 2.12 ;
        RECT  10.09 1.96 10.97 2.12 ;
        RECT  10.81 1.96 10.97 2.64 ;
        RECT  10.81 2.48 11.44 2.64 ;
        RECT  11.16 2.48 11.44 2.76 ;
        RECT  11.13 0.88 11.41 1.16 ;
        RECT  10.43 1.46 11.55 1.62 ;
        RECT  10.43 1.40 10.71 1.68 ;
        RECT  11.25 1.40 11.55 1.68 ;
        RECT  11.25 0.88 11.41 2.12 ;
        RECT  11.13 1.84 11.41 2.12 ;
    END
END DFFSSZSP2V1_0

MACRO DFFSSZSP1V1_0
    CLASS CORE ;
    FOREIGN DFFSSZSP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 23.49  LAYER ME1  ;
        ANTENNADIFFAREA 9.52  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.54  LAYER ME1  ;
        ANTENNAMAXAREACAR 43.69  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.73 1.46 12.34 1.74 ;
        RECT  11.61 1.90 11.89 2.18 ;
        RECT  11.73 0.96 11.89 2.18 ;
        RECT  11.61 0.96 11.89 1.24 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.52 1.40 9.94 1.68 ;
        END
    END SB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.24 1.40 3.54 1.76 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.20  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.83  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.81 1.19 2.25 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  0.91 0.81 1.19 1.09 ;
        END
    END D
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END SEL
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.87  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 12.90  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.06 1.46 2.34 1.74 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.81 2.23 2.25 ;
        RECT  1.95 0.81 2.23 1.09 ;
        END
    END TD
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 12.80 3.48 ;
        RECT  12.19 2.88 12.62 3.48 ;
        RECT  12.13 1.90 12.41 2.18 ;
        RECT  12.19 1.90 12.35 3.48 ;
        RECT  10.37 2.40 10.65 3.48 ;
        RECT  9.57 1.84 9.85 2.12 ;
        RECT  9.63 1.84 9.79 3.48 ;
        RECT  8.57 1.84 8.85 2.12 ;
        RECT  8.63 1.84 8.79 3.48 ;
        RECT  7.57 1.84 7.85 2.12 ;
        RECT  7.67 1.84 7.83 3.48 ;
        RECT  2.71 2.52 2.99 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 12.80 0.28 ;
        RECT  12.19 -0.28 12.62 0.32 ;
        RECT  12.13 0.96 12.41 1.24 ;
        RECT  12.19 -0.28 12.35 1.24 ;
        RECT  10.61 0.88 10.89 1.16 ;
        RECT  10.67 -0.28 10.83 1.16 ;
        RECT  9.13 -0.28 9.41 0.68 ;
        RECT  2.71 -0.28 2.99 0.68 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  1.55 1.97 1.71 2.57 ;
        RECT  1.55 2.41 2.37 2.57 ;
        RECT  2.09 2.41 2.37 2.69 ;
        RECT  3.47 0.96 3.86 1.24 ;
        RECT  3.70 1.46 4.02 1.74 ;
        RECT  3.70 0.96 3.86 2.20 ;
        RECT  3.47 1.92 3.86 2.20 ;
        RECT  4.07 0.44 4.35 0.72 ;
        RECT  3.15 0.56 4.35 0.72 ;
        RECT  3.15 0.56 3.31 1.12 ;
        RECT  2.43 0.96 3.31 1.12 ;
        RECT  2.43 0.96 2.71 1.24 ;
        RECT  2.55 0.96 2.71 2.20 ;
        RECT  2.43 1.92 2.71 2.20 ;
        RECT  2.43 2.04 3.31 2.20 ;
        RECT  3.15 2.04 3.31 2.64 ;
        RECT  3.15 2.48 4.25 2.64 ;
        RECT  3.97 2.48 4.25 2.76 ;
        RECT  5.59 0.76 5.91 1.04 ;
        RECT  5.59 0.76 5.75 2.00 ;
        RECT  5.25 1.84 6.29 2.00 ;
        RECT  5.25 1.84 5.53 2.12 ;
        RECT  6.01 1.84 6.29 2.12 ;
        RECT  6.15 0.76 6.43 1.04 ;
        RECT  6.27 0.76 6.43 1.36 ;
        RECT  7.11 1.08 7.39 1.36 ;
        RECT  6.27 1.20 7.39 1.36 ;
        RECT  6.53 1.20 6.69 2.12 ;
        RECT  6.53 1.84 6.81 2.12 ;
        RECT  4.63 0.86 4.91 1.14 ;
        RECT  4.07 0.98 4.91 1.14 ;
        RECT  4.07 0.96 4.35 1.24 ;
        RECT  4.29 0.98 4.45 2.12 ;
        RECT  4.41 1.84 4.57 2.44 ;
        RECT  4.41 2.28 7.51 2.44 ;
        RECT  7.23 2.28 7.51 2.56 ;
        RECT  6.67 0.76 7.95 0.92 ;
        RECT  6.67 0.76 6.95 1.04 ;
        RECT  7.67 0.76 7.95 1.16 ;
        RECT  7.67 0.76 7.83 1.68 ;
        RECT  8.71 1.40 8.99 1.68 ;
        RECT  7.25 1.52 8.99 1.68 ;
        RECT  8.01 1.52 8.17 2.12 ;
        RECT  7.25 1.52 7.41 2.12 ;
        RECT  7.05 1.84 7.41 2.12 ;
        RECT  8.01 1.84 8.37 2.12 ;
        RECT  5.27 0.44 8.87 0.60 ;
        RECT  8.71 0.44 8.87 1.04 ;
        RECT  8.71 0.88 9.37 1.04 ;
        RECT  5.27 0.44 5.43 1.14 ;
        RECT  9.09 0.88 9.37 1.16 ;
        RECT  5.15 0.86 5.31 1.46 ;
        RECT  4.93 1.30 5.31 1.46 ;
        RECT  9.15 0.88 9.31 2.12 ;
        RECT  4.93 1.30 5.09 2.12 ;
        RECT  4.81 1.84 5.09 2.12 ;
        RECT  9.09 1.84 9.37 2.12 ;
        RECT  9.71 0.88 9.99 1.16 ;
        RECT  9.71 1.00 10.26 1.16 ;
        RECT  10.10 1.00 10.26 2.12 ;
        RECT  10.09 1.84 10.37 2.12 ;
        RECT  10.09 1.96 10.97 2.12 ;
        RECT  10.81 1.96 10.97 2.64 ;
        RECT  10.81 2.48 11.44 2.64 ;
        RECT  11.16 2.48 11.44 2.76 ;
        RECT  11.13 0.88 11.41 1.16 ;
        RECT  10.43 1.46 11.55 1.62 ;
        RECT  10.43 1.40 10.71 1.68 ;
        RECT  11.25 1.40 11.55 1.68 ;
        RECT  11.25 0.88 11.41 2.12 ;
        RECT  11.13 1.84 11.41 2.12 ;
    END
END DFFSSZSP1V1_0

MACRO DFFSSSP8V1_0
    CLASS CORE ;
    FOREIGN DFFSSSP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.40 1.16 1.76 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.40 0.70 1.76 ;
        END
    END D
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.18 1.40 7.60 1.68 ;
        END
    END SB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 23.65  LAYER ME1  ;
        ANTENNADIFFAREA 11.24  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.98  LAYER ME1  ;
        ANTENNAMAXAREACAR 24.15  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.84 1.90 11.12 2.50 ;
        RECT  10.84 0.64 11.12 1.24 ;
        RECT  10.84 0.64 11.00 2.50 ;
        RECT  9.92 1.52 11.00 1.68 ;
        RECT  9.92 1.46 10.34 1.74 ;
        RECT  9.80 1.90 10.08 2.50 ;
        RECT  9.92 0.64 10.08 2.50 ;
        RECT  9.80 0.64 10.08 1.24 ;
        END
    END Q
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 12.00 3.48 ;
        RECT  11.42 2.88 11.82 3.48 ;
        RECT  11.36 1.90 11.64 2.50 ;
        RECT  11.42 1.90 11.58 3.48 ;
        RECT  10.32 1.90 10.60 2.50 ;
        RECT  10.38 1.90 10.54 3.48 ;
        RECT  9.28 1.90 9.56 2.50 ;
        RECT  9.34 1.90 9.50 3.48 ;
        RECT  8.04 2.40 8.32 3.48 ;
        RECT  7.24 1.84 7.52 2.12 ;
        RECT  7.30 1.84 7.46 3.48 ;
        RECT  6.24 1.84 6.52 2.12 ;
        RECT  6.30 1.84 6.46 3.48 ;
        RECT  5.24 1.84 5.52 2.12 ;
        RECT  5.34 1.84 5.50 3.48 ;
        RECT  0.38 2.48 0.66 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 12.00 0.28 ;
        RECT  11.42 -0.28 11.82 0.32 ;
        RECT  11.36 0.64 11.64 1.24 ;
        RECT  11.42 -0.28 11.58 1.24 ;
        RECT  10.32 0.64 10.60 1.24 ;
        RECT  10.38 -0.28 10.54 1.24 ;
        RECT  9.28 0.64 9.56 1.24 ;
        RECT  9.34 -0.28 9.50 1.24 ;
        RECT  8.28 0.88 8.56 1.16 ;
        RECT  8.34 -0.28 8.50 1.16 ;
        RECT  6.80 -0.28 7.08 0.68 ;
        RECT  0.38 -0.28 0.66 0.68 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  1.14 0.96 1.48 1.24 ;
        RECT  1.32 1.46 1.64 1.74 ;
        RECT  1.32 0.96 1.48 2.20 ;
        RECT  1.14 1.92 1.48 2.20 ;
        RECT  1.74 0.44 2.02 0.72 ;
        RECT  0.82 0.56 2.02 0.72 ;
        RECT  0.82 0.56 0.98 1.12 ;
        RECT  0.08 0.96 0.98 1.12 ;
        RECT  0.08 0.96 0.38 1.24 ;
        RECT  0.08 0.96 0.24 2.20 ;
        RECT  0.08 1.92 0.38 2.20 ;
        RECT  0.08 2.04 0.98 2.20 ;
        RECT  0.82 2.04 0.98 2.64 ;
        RECT  0.82 2.48 1.92 2.64 ;
        RECT  1.64 2.48 1.92 2.76 ;
        RECT  3.26 0.76 3.58 1.04 ;
        RECT  3.26 0.76 3.42 2.00 ;
        RECT  2.92 1.84 3.96 2.00 ;
        RECT  2.92 1.84 3.20 2.12 ;
        RECT  3.68 1.84 3.96 2.12 ;
        RECT  3.82 0.76 4.10 1.04 ;
        RECT  3.94 0.76 4.10 1.36 ;
        RECT  4.78 1.08 5.06 1.36 ;
        RECT  3.94 1.20 5.06 1.36 ;
        RECT  4.20 1.20 4.36 2.12 ;
        RECT  4.20 1.84 4.48 2.12 ;
        RECT  2.30 0.86 2.58 1.14 ;
        RECT  1.74 0.98 2.58 1.14 ;
        RECT  1.74 0.96 2.02 1.24 ;
        RECT  1.96 0.98 2.12 2.12 ;
        RECT  2.08 1.84 2.24 2.44 ;
        RECT  2.08 2.28 5.18 2.44 ;
        RECT  4.90 2.28 5.18 2.56 ;
        RECT  4.34 0.76 5.62 0.92 ;
        RECT  4.34 0.76 4.62 1.04 ;
        RECT  5.34 0.76 5.62 1.16 ;
        RECT  5.34 0.76 5.50 1.68 ;
        RECT  6.38 1.40 6.66 1.68 ;
        RECT  4.92 1.52 6.66 1.68 ;
        RECT  5.68 1.52 5.84 2.12 ;
        RECT  4.92 1.52 5.08 2.12 ;
        RECT  4.72 1.84 5.08 2.12 ;
        RECT  5.68 1.84 6.04 2.12 ;
        RECT  2.94 0.44 6.54 0.60 ;
        RECT  6.38 0.44 6.54 1.04 ;
        RECT  6.38 0.88 7.04 1.04 ;
        RECT  2.94 0.44 3.10 1.14 ;
        RECT  6.76 0.88 7.04 1.16 ;
        RECT  2.82 0.86 2.98 1.46 ;
        RECT  2.60 1.30 2.98 1.46 ;
        RECT  6.82 0.88 6.98 2.12 ;
        RECT  2.60 1.30 2.76 2.12 ;
        RECT  2.48 1.84 2.76 2.12 ;
        RECT  6.76 1.84 7.04 2.12 ;
        RECT  7.38 0.88 7.66 1.16 ;
        RECT  7.38 1.00 7.92 1.16 ;
        RECT  7.76 1.00 7.92 2.12 ;
        RECT  7.76 1.84 8.04 2.12 ;
        RECT  7.76 1.96 8.64 2.12 ;
        RECT  8.48 1.96 8.64 2.64 ;
        RECT  8.48 2.48 9.11 2.64 ;
        RECT  8.83 2.48 9.11 2.76 ;
        RECT  8.80 0.88 9.08 1.16 ;
        RECT  8.10 1.46 9.22 1.62 ;
        RECT  8.10 1.40 8.38 1.68 ;
        RECT  8.92 1.40 9.22 1.68 ;
        RECT  8.92 0.88 9.08 2.12 ;
        RECT  8.80 1.84 9.08 2.12 ;
    END
END DFFSSSP8V1_0

MACRO DFFSSSP4V1_0
    CLASS CORE ;
    FOREIGN DFFSSSP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 21.31  LAYER ME1  ;
        ANTENNADIFFAREA 9.41  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.69  LAYER ME1  ;
        ANTENNAMAXAREACAR 30.83  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.92 1.46 10.34 1.74 ;
        RECT  9.80 1.90 10.08 2.50 ;
        RECT  9.92 0.64 10.08 2.50 ;
        RECT  9.80 0.64 10.08 1.24 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.18 1.40 7.60 1.68 ;
        END
    END SB
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.40 0.70 1.76 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.40 1.16 1.76 ;
        END
    END CK
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 10.80 0.28 ;
        RECT  10.34 -0.28 10.62 0.32 ;
        RECT  10.32 0.64 10.60 1.24 ;
        RECT  10.38 -0.28 10.54 1.24 ;
        RECT  9.28 0.64 9.56 1.24 ;
        RECT  9.34 -0.28 9.50 1.24 ;
        RECT  8.28 0.88 8.56 1.16 ;
        RECT  8.34 -0.28 8.50 1.16 ;
        RECT  6.80 -0.28 7.08 0.68 ;
        RECT  0.38 -0.28 0.66 0.68 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 10.80 3.48 ;
        RECT  10.34 2.88 10.62 3.48 ;
        RECT  10.32 1.90 10.60 2.50 ;
        RECT  10.38 1.90 10.54 3.48 ;
        RECT  9.28 1.90 9.56 2.50 ;
        RECT  9.34 1.90 9.50 3.48 ;
        RECT  8.04 2.40 8.32 3.48 ;
        RECT  7.24 1.84 7.52 2.12 ;
        RECT  7.30 1.84 7.46 3.48 ;
        RECT  6.24 1.84 6.52 2.12 ;
        RECT  6.30 1.84 6.46 3.48 ;
        RECT  5.24 1.84 5.52 2.12 ;
        RECT  5.34 1.84 5.50 3.48 ;
        RECT  0.38 2.48 0.66 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  1.14 0.96 1.48 1.24 ;
        RECT  1.32 1.46 1.64 1.74 ;
        RECT  1.32 0.96 1.48 2.20 ;
        RECT  1.14 1.92 1.48 2.20 ;
        RECT  1.74 0.44 2.02 0.72 ;
        RECT  0.82 0.56 2.02 0.72 ;
        RECT  0.82 0.56 0.98 1.12 ;
        RECT  0.08 0.96 0.98 1.12 ;
        RECT  0.08 0.96 0.38 1.24 ;
        RECT  0.08 0.96 0.24 2.20 ;
        RECT  0.08 1.92 0.38 2.20 ;
        RECT  0.08 2.04 0.98 2.20 ;
        RECT  0.82 2.04 0.98 2.64 ;
        RECT  0.82 2.48 1.92 2.64 ;
        RECT  1.64 2.48 1.92 2.76 ;
        RECT  3.26 0.76 3.58 1.04 ;
        RECT  3.26 0.76 3.42 2.00 ;
        RECT  2.92 1.84 3.96 2.00 ;
        RECT  2.92 1.84 3.20 2.12 ;
        RECT  3.68 1.84 3.96 2.12 ;
        RECT  3.82 0.76 4.10 1.04 ;
        RECT  3.94 0.76 4.10 1.36 ;
        RECT  4.78 1.08 5.06 1.36 ;
        RECT  3.94 1.20 5.06 1.36 ;
        RECT  4.20 1.20 4.36 2.12 ;
        RECT  4.20 1.84 4.48 2.12 ;
        RECT  2.30 0.86 2.58 1.14 ;
        RECT  1.74 0.98 2.58 1.14 ;
        RECT  1.74 0.96 2.02 1.24 ;
        RECT  1.96 0.98 2.12 2.12 ;
        RECT  2.08 1.84 2.24 2.44 ;
        RECT  2.08 2.28 5.18 2.44 ;
        RECT  4.90 2.28 5.18 2.56 ;
        RECT  4.34 0.76 5.62 0.92 ;
        RECT  4.34 0.76 4.62 1.04 ;
        RECT  5.34 0.76 5.62 1.16 ;
        RECT  5.34 0.76 5.50 1.68 ;
        RECT  6.38 1.40 6.66 1.68 ;
        RECT  4.92 1.52 6.66 1.68 ;
        RECT  5.68 1.52 5.84 2.12 ;
        RECT  4.92 1.52 5.08 2.12 ;
        RECT  4.72 1.84 5.08 2.12 ;
        RECT  5.68 1.84 6.04 2.12 ;
        RECT  2.94 0.44 6.54 0.60 ;
        RECT  6.38 0.44 6.54 1.04 ;
        RECT  6.38 0.88 7.04 1.04 ;
        RECT  2.94 0.44 3.10 1.14 ;
        RECT  6.76 0.88 7.04 1.16 ;
        RECT  2.82 0.86 2.98 1.46 ;
        RECT  2.60 1.30 2.98 1.46 ;
        RECT  6.82 0.88 6.98 2.12 ;
        RECT  2.60 1.30 2.76 2.12 ;
        RECT  2.48 1.84 2.76 2.12 ;
        RECT  6.76 1.84 7.04 2.12 ;
        RECT  7.38 0.88 7.66 1.16 ;
        RECT  7.38 1.00 7.92 1.16 ;
        RECT  7.76 1.00 7.92 2.12 ;
        RECT  7.76 1.84 8.04 2.12 ;
        RECT  7.76 1.96 8.64 2.12 ;
        RECT  8.48 1.96 8.64 2.64 ;
        RECT  8.48 2.48 9.11 2.64 ;
        RECT  8.83 2.48 9.11 2.76 ;
        RECT  8.80 0.88 9.08 1.16 ;
        RECT  8.10 1.46 9.22 1.62 ;
        RECT  8.10 1.40 8.38 1.68 ;
        RECT  8.92 1.40 9.22 1.68 ;
        RECT  8.92 0.88 9.08 2.12 ;
        RECT  8.80 1.84 9.08 2.12 ;
    END
END DFFSSSP4V1_0

MACRO DFFSSSP2V1_0
    CLASS CORE ;
    FOREIGN DFFSSSP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.40 1.16 1.76 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.40 0.70 1.76 ;
        END
    END D
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.18 1.40 7.60 1.68 ;
        END
    END SB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 20.44  LAYER ME1  ;
        ANTENNADIFFAREA 8.80  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.55  LAYER ME1  ;
        ANTENNAMAXAREACAR 37.35  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.40 1.46 9.94 1.74 ;
        RECT  9.28 1.90 9.56 2.50 ;
        RECT  9.40 0.64 9.56 2.50 ;
        RECT  9.28 0.64 9.56 1.24 ;
        END
    END Q
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 10.40 3.48 ;
        RECT  9.86 2.88 10.22 3.48 ;
        RECT  9.80 1.90 10.08 2.50 ;
        RECT  9.86 1.90 10.02 3.48 ;
        RECT  8.04 2.40 8.32 3.48 ;
        RECT  7.24 1.84 7.52 2.12 ;
        RECT  7.30 1.84 7.46 3.48 ;
        RECT  6.24 1.84 6.52 2.12 ;
        RECT  6.30 1.84 6.46 3.48 ;
        RECT  5.24 1.84 5.52 2.12 ;
        RECT  5.34 1.84 5.50 3.48 ;
        RECT  0.38 2.48 0.66 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 10.40 0.28 ;
        RECT  9.86 -0.28 10.22 0.32 ;
        RECT  9.80 0.64 10.08 1.24 ;
        RECT  9.86 -0.28 10.02 1.24 ;
        RECT  8.28 0.88 8.56 1.16 ;
        RECT  8.34 -0.28 8.50 1.16 ;
        RECT  6.80 -0.28 7.08 0.68 ;
        RECT  0.38 -0.28 0.66 0.68 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  1.14 0.96 1.48 1.24 ;
        RECT  1.32 1.46 1.64 1.74 ;
        RECT  1.32 0.96 1.48 2.20 ;
        RECT  1.14 1.92 1.48 2.20 ;
        RECT  1.74 0.44 2.02 0.72 ;
        RECT  0.82 0.56 2.02 0.72 ;
        RECT  0.82 0.56 0.98 1.12 ;
        RECT  0.08 0.96 0.98 1.12 ;
        RECT  0.08 0.96 0.38 1.24 ;
        RECT  0.08 0.96 0.24 2.20 ;
        RECT  0.08 1.92 0.38 2.20 ;
        RECT  0.08 2.04 0.98 2.20 ;
        RECT  0.82 2.04 0.98 2.64 ;
        RECT  0.82 2.48 1.92 2.64 ;
        RECT  1.64 2.48 1.92 2.76 ;
        RECT  3.26 0.76 3.58 1.04 ;
        RECT  3.26 0.76 3.42 2.00 ;
        RECT  2.92 1.84 3.96 2.00 ;
        RECT  2.92 1.84 3.20 2.12 ;
        RECT  3.68 1.84 3.96 2.12 ;
        RECT  3.82 0.76 4.10 1.04 ;
        RECT  3.94 0.76 4.10 1.36 ;
        RECT  4.78 1.08 5.06 1.36 ;
        RECT  3.94 1.20 5.06 1.36 ;
        RECT  4.20 1.20 4.36 2.12 ;
        RECT  4.20 1.84 4.48 2.12 ;
        RECT  2.30 0.86 2.58 1.14 ;
        RECT  1.74 0.98 2.58 1.14 ;
        RECT  1.74 0.96 2.02 1.24 ;
        RECT  1.96 0.98 2.12 2.12 ;
        RECT  2.08 1.84 2.24 2.44 ;
        RECT  2.08 2.28 5.18 2.44 ;
        RECT  4.90 2.28 5.18 2.56 ;
        RECT  4.34 0.76 5.62 0.92 ;
        RECT  4.34 0.76 4.62 1.04 ;
        RECT  5.34 0.76 5.62 1.16 ;
        RECT  5.34 0.76 5.50 1.68 ;
        RECT  6.38 1.40 6.66 1.68 ;
        RECT  4.92 1.52 6.66 1.68 ;
        RECT  5.68 1.52 5.84 2.12 ;
        RECT  4.92 1.52 5.08 2.12 ;
        RECT  4.72 1.84 5.08 2.12 ;
        RECT  5.68 1.84 6.04 2.12 ;
        RECT  2.94 0.44 6.54 0.60 ;
        RECT  6.38 0.44 6.54 1.04 ;
        RECT  6.38 0.88 7.04 1.04 ;
        RECT  2.94 0.44 3.10 1.14 ;
        RECT  6.76 0.88 7.04 1.16 ;
        RECT  2.82 0.86 2.98 1.46 ;
        RECT  2.60 1.30 2.98 1.46 ;
        RECT  6.82 0.88 6.98 2.12 ;
        RECT  2.60 1.30 2.76 2.12 ;
        RECT  2.48 1.84 2.76 2.12 ;
        RECT  6.76 1.84 7.04 2.12 ;
        RECT  7.38 0.88 7.66 1.16 ;
        RECT  7.38 1.00 7.92 1.16 ;
        RECT  7.76 1.00 7.92 2.12 ;
        RECT  7.76 1.84 8.04 2.12 ;
        RECT  7.76 1.96 8.64 2.12 ;
        RECT  8.48 1.96 8.64 2.64 ;
        RECT  8.48 2.48 9.11 2.64 ;
        RECT  8.83 2.48 9.11 2.76 ;
        RECT  8.80 0.88 9.08 1.16 ;
        RECT  8.10 1.46 9.22 1.62 ;
        RECT  8.10 1.40 8.38 1.68 ;
        RECT  8.92 1.40 9.22 1.68 ;
        RECT  8.92 0.88 9.08 2.12 ;
        RECT  8.80 1.84 9.08 2.12 ;
    END
END DFFSSSP2V1_0

MACRO DFFSSSP1V1_0
    CLASS CORE ;
    FOREIGN DFFSSSP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.40 0.70 1.76 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.40 1.16 1.76 ;
        END
    END CK
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.18 1.40 7.60 1.68 ;
        END
    END SB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 20.18  LAYER ME1  ;
        ANTENNADIFFAREA 8.37  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.47  LAYER ME1  ;
        ANTENNAMAXAREACAR 42.91  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.40 1.46 9.94 1.74 ;
        RECT  9.28 1.90 9.56 2.18 ;
        RECT  9.40 0.96 9.56 2.18 ;
        RECT  9.28 0.96 9.56 1.24 ;
        END
    END Q
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 10.40 0.28 ;
        RECT  9.86 -0.28 10.22 0.32 ;
        RECT  9.80 0.96 10.08 1.24 ;
        RECT  9.86 -0.28 10.02 1.24 ;
        RECT  8.28 0.88 8.56 1.16 ;
        RECT  8.34 -0.28 8.50 1.16 ;
        RECT  6.80 -0.28 7.08 0.68 ;
        RECT  0.38 -0.28 0.66 0.68 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 10.40 3.48 ;
        RECT  9.86 2.88 10.22 3.48 ;
        RECT  9.80 1.90 10.08 2.18 ;
        RECT  9.86 1.90 10.02 3.48 ;
        RECT  8.04 2.40 8.32 3.48 ;
        RECT  7.24 1.84 7.52 2.12 ;
        RECT  7.30 1.84 7.46 3.48 ;
        RECT  6.24 1.84 6.52 2.12 ;
        RECT  6.30 1.84 6.46 3.48 ;
        RECT  5.24 1.84 5.52 2.12 ;
        RECT  5.34 1.84 5.50 3.48 ;
        RECT  0.38 2.48 0.66 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  1.14 0.96 1.48 1.24 ;
        RECT  1.32 1.46 1.64 1.74 ;
        RECT  1.32 0.96 1.48 2.20 ;
        RECT  1.14 1.92 1.48 2.20 ;
        RECT  1.74 0.44 2.02 0.72 ;
        RECT  0.82 0.56 2.02 0.72 ;
        RECT  0.82 0.56 0.98 1.12 ;
        RECT  0.08 0.96 0.98 1.12 ;
        RECT  0.08 0.96 0.38 1.24 ;
        RECT  0.08 0.96 0.24 2.20 ;
        RECT  0.08 1.92 0.38 2.20 ;
        RECT  0.08 2.04 0.98 2.20 ;
        RECT  0.82 2.04 0.98 2.64 ;
        RECT  0.82 2.48 1.92 2.64 ;
        RECT  1.64 2.48 1.92 2.76 ;
        RECT  3.26 0.76 3.58 1.04 ;
        RECT  3.26 0.76 3.42 2.00 ;
        RECT  2.92 1.84 3.96 2.00 ;
        RECT  2.92 1.84 3.20 2.12 ;
        RECT  3.68 1.84 3.96 2.12 ;
        RECT  3.82 0.76 4.10 1.04 ;
        RECT  3.94 0.76 4.10 1.36 ;
        RECT  4.78 1.08 5.06 1.36 ;
        RECT  3.94 1.20 5.06 1.36 ;
        RECT  4.20 1.20 4.36 2.12 ;
        RECT  4.20 1.84 4.48 2.12 ;
        RECT  2.30 0.86 2.58 1.14 ;
        RECT  1.74 0.98 2.58 1.14 ;
        RECT  1.74 0.96 2.02 1.24 ;
        RECT  1.96 0.98 2.12 2.12 ;
        RECT  2.08 1.84 2.24 2.44 ;
        RECT  2.08 2.28 5.18 2.44 ;
        RECT  4.90 2.28 5.18 2.56 ;
        RECT  4.34 0.76 5.62 0.92 ;
        RECT  4.34 0.76 4.62 1.04 ;
        RECT  5.34 0.76 5.62 1.16 ;
        RECT  5.34 0.76 5.50 1.68 ;
        RECT  6.38 1.40 6.66 1.68 ;
        RECT  4.92 1.52 6.66 1.68 ;
        RECT  5.68 1.52 5.84 2.12 ;
        RECT  4.92 1.52 5.08 2.12 ;
        RECT  4.72 1.84 5.08 2.12 ;
        RECT  5.68 1.84 6.04 2.12 ;
        RECT  2.94 0.44 6.54 0.60 ;
        RECT  6.38 0.44 6.54 1.04 ;
        RECT  6.38 0.88 7.04 1.04 ;
        RECT  2.94 0.44 3.10 1.14 ;
        RECT  6.76 0.88 7.04 1.16 ;
        RECT  2.82 0.86 2.98 1.46 ;
        RECT  2.60 1.30 2.98 1.46 ;
        RECT  6.82 0.88 6.98 2.12 ;
        RECT  2.60 1.30 2.76 2.12 ;
        RECT  2.48 1.84 2.76 2.12 ;
        RECT  6.76 1.84 7.04 2.12 ;
        RECT  7.38 0.88 7.66 1.16 ;
        RECT  7.38 1.00 7.92 1.16 ;
        RECT  7.76 1.00 7.92 2.12 ;
        RECT  7.76 1.84 8.04 2.12 ;
        RECT  7.76 1.96 8.64 2.12 ;
        RECT  8.48 1.96 8.64 2.64 ;
        RECT  8.48 2.48 9.11 2.64 ;
        RECT  8.83 2.48 9.11 2.76 ;
        RECT  8.80 0.88 9.08 1.16 ;
        RECT  8.10 1.46 9.22 1.62 ;
        RECT  8.10 1.40 8.38 1.68 ;
        RECT  8.92 1.40 9.22 1.68 ;
        RECT  8.92 0.88 9.08 2.12 ;
        RECT  8.80 1.84 9.08 2.12 ;
    END
END DFFSSSP1V1_0

MACRO DFFSSP8V1_1
    CLASS CORE ;
    FOREIGN DFFSSP8V1_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 17.91  LAYER ME1  ;
        ANTENNADIFFAREA 8.84  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.98  LAYER ME1  ;
        ANTENNAMAXAREACAR 18.30  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.64 1.84 8.92 2.12 ;
        RECT  8.64 0.96 8.92 1.24 ;
        RECT  8.64 0.96 8.80 2.12 ;
        RECT  7.66 1.52 8.80 1.68 ;
        RECT  7.66 1.46 7.92 1.74 ;
        RECT  7.60 1.84 7.88 2.12 ;
        RECT  7.66 0.96 7.88 2.12 ;
        RECT  7.60 0.96 7.88 1.24 ;
        END
    END Q
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.88 1.39 1.16 1.81 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.39 0.72 1.81 ;
        END
    END D
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 9.60 0.28 ;
        RECT  9.16 0.64 9.44 0.92 ;
        RECT  9.14 -0.28 9.42 0.32 ;
        RECT  9.22 -0.28 9.38 0.92 ;
        RECT  8.12 0.64 8.40 0.92 ;
        RECT  8.18 -0.28 8.34 0.92 ;
        RECT  7.08 0.64 7.36 0.92 ;
        RECT  7.14 -0.28 7.30 0.92 ;
        RECT  6.08 0.96 6.36 1.24 ;
        RECT  6.18 -0.28 6.34 1.24 ;
        RECT  3.36 0.72 3.64 1.00 ;
        RECT  3.42 -0.28 3.58 1.00 ;
        RECT  0.62 0.68 0.90 0.96 ;
        RECT  0.68 -0.28 0.84 0.96 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 9.60 3.48 ;
        RECT  9.16 2.16 9.44 2.44 ;
        RECT  9.14 2.88 9.42 3.48 ;
        RECT  9.22 2.16 9.38 3.48 ;
        RECT  8.12 2.16 8.40 2.44 ;
        RECT  8.18 2.16 8.34 3.48 ;
        RECT  7.08 2.16 7.36 2.44 ;
        RECT  7.14 2.16 7.30 3.48 ;
        RECT  6.08 2.62 6.36 3.48 ;
        RECT  3.48 1.92 3.76 2.20 ;
        RECT  3.54 1.92 3.70 3.48 ;
        RECT  0.38 2.62 0.66 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  1.14 0.68 1.48 0.96 ;
        RECT  1.32 1.22 1.64 1.50 ;
        RECT  1.32 0.68 1.48 2.25 ;
        RECT  1.14 1.97 1.48 2.25 ;
        RECT  0.08 0.68 0.38 0.96 ;
        RECT  1.68 0.72 1.96 1.00 ;
        RECT  0.08 0.68 0.24 2.25 ;
        RECT  0.08 1.97 0.38 2.25 ;
        RECT  1.80 0.72 1.96 2.20 ;
        RECT  0.08 2.09 0.98 2.25 ;
        RECT  0.82 2.09 0.98 2.57 ;
        RECT  1.68 1.92 1.84 2.57 ;
        RECT  0.82 2.41 1.84 2.57 ;
        RECT  2.76 0.72 3.07 1.00 ;
        RECT  2.76 0.72 2.92 2.20 ;
        RECT  2.72 1.92 3.00 2.20 ;
        RECT  2.20 0.72 2.48 1.00 ;
        RECT  3.56 1.48 3.84 1.76 ;
        RECT  3.16 1.60 3.84 1.76 ;
        RECT  2.26 0.72 2.42 2.20 ;
        RECT  2.20 1.92 2.48 2.20 ;
        RECT  2.32 1.92 2.48 2.52 ;
        RECT  3.16 1.60 3.32 2.52 ;
        RECT  2.32 2.36 3.32 2.52 ;
        RECT  3.88 0.72 4.16 1.00 ;
        RECT  3.08 1.16 4.16 1.32 ;
        RECT  3.08 1.16 3.36 1.44 ;
        RECT  4.00 0.72 4.16 2.20 ;
        RECT  4.00 1.92 4.28 2.20 ;
        RECT  4.56 0.44 6.02 0.60 ;
        RECT  5.74 0.44 6.02 0.80 ;
        RECT  4.44 0.76 4.72 1.04 ;
        RECT  4.56 0.44 4.72 2.20 ;
        RECT  4.52 1.92 4.80 2.20 ;
        RECT  5.56 0.96 5.84 1.24 ;
        RECT  5.56 1.46 6.56 1.62 ;
        RECT  6.28 1.40 6.56 1.68 ;
        RECT  5.56 0.96 5.72 2.12 ;
        RECT  5.56 1.84 5.84 2.12 ;
        RECT  4.96 0.76 5.24 1.04 ;
        RECT  6.60 0.96 6.88 1.24 ;
        RECT  6.60 1.84 6.88 2.12 ;
        RECT  5.08 0.76 5.24 2.20 ;
        RECT  5.04 1.92 5.32 2.20 ;
        RECT  5.16 1.92 5.32 2.44 ;
        RECT  6.72 0.96 6.88 2.44 ;
        RECT  5.16 2.28 6.88 2.44 ;
    END
END DFFSSP8V1_1

MACRO DFFSSP8V1_0
    CLASS CORE ;
    FOREIGN DFFSSP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 17.86  LAYER ME1  ;
        ANTENNADIFFAREA 9.26  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.23  LAYER ME1  ;
        ANTENNAMAXAREACAR 14.48  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.58 1.92 8.86 2.20 ;
        RECT  8.58 0.96 8.86 1.24 ;
        RECT  8.58 0.96 8.74 2.20 ;
        RECT  7.72 1.52 8.74 1.68 ;
        RECT  7.54 1.92 7.88 2.20 ;
        RECT  7.72 0.96 7.88 2.20 ;
        RECT  7.54 0.96 7.88 1.24 ;
        END
    END Q
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.40 0.82 1.68 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.72 1.40 2.14 1.68 ;
        END
    END D
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 9.60 0.28 ;
        RECT  9.14 -0.28 9.42 0.32 ;
        RECT  9.10 0.62 9.38 0.90 ;
        RECT  9.16 -0.28 9.32 0.90 ;
        RECT  8.06 0.62 8.34 0.90 ;
        RECT  8.12 -0.28 8.28 0.90 ;
        RECT  7.02 0.62 7.30 0.90 ;
        RECT  7.08 -0.28 7.24 0.90 ;
        RECT  5.90 0.72 6.18 1.00 ;
        RECT  5.96 -0.28 6.12 1.00 ;
        RECT  3.82 0.72 4.10 1.00 ;
        RECT  3.88 -0.28 4.04 1.00 ;
        RECT  1.74 0.72 2.02 1.00 ;
        RECT  1.80 -0.28 1.96 1.00 ;
        RECT  0.62 0.52 0.90 0.80 ;
        RECT  0.68 -0.28 0.84 0.80 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 9.60 3.48 ;
        RECT  9.14 2.88 9.42 3.48 ;
        RECT  9.10 2.26 9.38 2.54 ;
        RECT  9.16 2.26 9.32 3.48 ;
        RECT  8.06 2.26 8.34 2.54 ;
        RECT  8.12 2.26 8.28 3.48 ;
        RECT  7.02 2.26 7.30 2.54 ;
        RECT  7.08 2.26 7.24 3.48 ;
        RECT  6.14 2.52 6.42 3.48 ;
        RECT  4.06 2.52 4.34 3.48 ;
        RECT  1.74 1.92 2.02 2.20 ;
        RECT  1.80 1.92 1.96 3.48 ;
        RECT  0.62 1.84 0.90 2.12 ;
        RECT  0.68 1.84 0.84 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.08 0.52 0.38 0.80 ;
        RECT  0.08 1.01 1.10 1.17 ;
        RECT  0.82 0.96 1.10 1.24 ;
        RECT  0.08 0.52 0.24 2.12 ;
        RECT  0.08 1.84 0.38 2.12 ;
        RECT  1.14 0.52 1.42 0.80 ;
        RECT  1.26 1.40 1.56 1.68 ;
        RECT  1.26 0.52 1.42 2.12 ;
        RECT  1.14 1.84 1.42 2.12 ;
        RECT  2.26 0.72 2.54 1.00 ;
        RECT  2.32 0.72 2.48 2.20 ;
        RECT  2.26 1.92 2.54 2.20 ;
        RECT  3.24 0.72 3.58 1.00 ;
        RECT  3.24 0.72 3.40 2.20 ;
        RECT  3.24 1.92 3.58 2.20 ;
        RECT  2.78 0.72 3.06 1.00 ;
        RECT  4.04 1.48 4.32 1.76 ;
        RECT  3.74 1.60 4.32 1.76 ;
        RECT  2.84 0.72 3.00 2.20 ;
        RECT  2.78 1.92 3.06 2.20 ;
        RECT  2.90 1.92 3.06 2.52 ;
        RECT  3.74 1.60 3.90 2.52 ;
        RECT  2.90 2.36 3.90 2.52 ;
        RECT  4.34 0.72 4.64 1.00 ;
        RECT  3.56 1.16 4.64 1.32 ;
        RECT  3.56 1.16 3.84 1.44 ;
        RECT  4.48 0.72 4.64 2.20 ;
        RECT  4.34 1.92 4.64 2.20 ;
        RECT  5.32 0.72 5.66 1.00 ;
        RECT  5.32 0.72 5.48 2.20 ;
        RECT  5.32 1.92 5.66 2.20 ;
        RECT  4.86 0.72 5.14 1.00 ;
        RECT  6.12 1.48 6.40 1.76 ;
        RECT  5.82 1.60 6.40 1.76 ;
        RECT  4.92 0.72 5.08 2.20 ;
        RECT  4.86 1.92 5.14 2.20 ;
        RECT  4.98 1.92 5.14 2.52 ;
        RECT  5.82 1.60 5.98 2.52 ;
        RECT  4.98 2.36 5.98 2.52 ;
        RECT  6.42 0.72 6.72 1.00 ;
        RECT  5.64 1.16 6.72 1.32 ;
        RECT  5.64 1.16 5.92 1.44 ;
        RECT  6.56 1.54 7.48 1.70 ;
        RECT  7.20 1.48 7.48 1.76 ;
        RECT  6.56 0.72 6.72 2.20 ;
        RECT  6.42 1.92 6.72 2.20 ;
    END
END DFFSSP8V1_0

MACRO DFFSSP4V1_1
    CLASS CORE ;
    FOREIGN DFFSSP4V1_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.39 0.72 1.81 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.88 1.39 1.16 1.81 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 16.07  LAYER ME1  ;
        ANTENNADIFFAREA 7.42  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.69  LAYER ME1  ;
        ANTENNAMAXAREACAR 23.25  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.66 1.46 7.92 1.74 ;
        RECT  7.60 1.84 7.88 2.12 ;
        RECT  7.66 0.96 7.88 2.12 ;
        RECT  7.60 0.96 7.88 1.24 ;
        END
    END Q
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 8.80 3.48 ;
        RECT  8.18 2.88 8.62 3.48 ;
        RECT  8.12 2.16 8.40 2.44 ;
        RECT  8.18 2.16 8.34 3.48 ;
        RECT  7.08 2.16 7.36 2.44 ;
        RECT  7.14 2.16 7.30 3.48 ;
        RECT  6.08 2.62 6.36 3.48 ;
        RECT  3.48 1.92 3.76 2.20 ;
        RECT  3.54 1.92 3.70 3.48 ;
        RECT  0.38 2.62 0.66 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 8.80 0.28 ;
        RECT  8.18 -0.28 8.62 0.32 ;
        RECT  8.12 0.64 8.40 0.92 ;
        RECT  8.18 -0.28 8.34 0.92 ;
        RECT  7.08 0.64 7.36 0.92 ;
        RECT  7.14 -0.28 7.30 0.92 ;
        RECT  6.08 0.96 6.36 1.24 ;
        RECT  6.18 -0.28 6.34 1.24 ;
        RECT  3.36 0.72 3.64 1.00 ;
        RECT  3.42 -0.28 3.58 1.00 ;
        RECT  0.62 0.68 0.90 0.96 ;
        RECT  0.68 -0.28 0.84 0.96 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  1.14 0.68 1.48 0.96 ;
        RECT  1.32 1.22 1.64 1.50 ;
        RECT  1.32 0.68 1.48 2.25 ;
        RECT  1.14 1.97 1.48 2.25 ;
        RECT  0.08 0.68 0.38 0.96 ;
        RECT  1.68 0.72 1.96 1.00 ;
        RECT  0.08 0.68 0.24 2.25 ;
        RECT  0.08 1.97 0.38 2.25 ;
        RECT  1.80 0.72 1.96 2.20 ;
        RECT  0.08 2.09 0.98 2.25 ;
        RECT  0.82 2.09 0.98 2.57 ;
        RECT  1.68 1.92 1.84 2.57 ;
        RECT  0.82 2.41 1.84 2.57 ;
        RECT  2.76 0.72 3.07 1.00 ;
        RECT  2.76 0.72 2.92 2.20 ;
        RECT  2.72 1.92 3.00 2.20 ;
        RECT  2.20 0.72 2.48 1.00 ;
        RECT  3.56 1.48 3.84 1.76 ;
        RECT  3.16 1.60 3.84 1.76 ;
        RECT  2.26 0.72 2.42 2.20 ;
        RECT  2.20 1.92 2.48 2.20 ;
        RECT  2.32 1.92 2.48 2.52 ;
        RECT  3.16 1.60 3.32 2.52 ;
        RECT  2.32 2.36 3.32 2.52 ;
        RECT  3.88 0.72 4.16 1.00 ;
        RECT  3.08 1.16 4.16 1.32 ;
        RECT  3.08 1.16 3.36 1.44 ;
        RECT  4.00 0.72 4.16 2.20 ;
        RECT  4.00 1.92 4.28 2.20 ;
        RECT  4.56 0.44 6.02 0.60 ;
        RECT  5.74 0.44 6.02 0.80 ;
        RECT  4.44 0.76 4.72 1.04 ;
        RECT  4.56 0.44 4.72 2.20 ;
        RECT  4.52 1.92 4.80 2.20 ;
        RECT  5.56 0.96 5.84 1.24 ;
        RECT  5.56 1.46 6.56 1.62 ;
        RECT  6.28 1.40 6.56 1.68 ;
        RECT  5.56 0.96 5.72 2.12 ;
        RECT  5.56 1.84 5.84 2.12 ;
        RECT  4.96 0.76 5.24 1.04 ;
        RECT  6.60 0.96 6.88 1.24 ;
        RECT  6.60 1.84 6.88 2.12 ;
        RECT  5.08 0.76 5.24 2.20 ;
        RECT  5.04 1.92 5.32 2.20 ;
        RECT  5.16 1.92 5.32 2.44 ;
        RECT  6.72 0.96 6.88 2.44 ;
        RECT  5.16 2.28 6.88 2.44 ;
    END
END DFFSSP4V1_1

MACRO DFFSSP4V1_0
    CLASS CORE ;
    FOREIGN DFFSSP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.72 1.40 2.14 1.68 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.40 0.82 1.68 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 16.01  LAYER ME1  ;
        ANTENNADIFFAREA 7.89  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.96  LAYER ME1  ;
        ANTENNAMAXAREACAR 16.76  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.54 1.92 7.88 2.20 ;
        RECT  7.72 0.96 7.88 2.20 ;
        RECT  7.54 0.96 7.88 1.24 ;
        END
    END Q
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 8.80 3.48 ;
        RECT  8.12 2.88 8.62 3.48 ;
        RECT  8.06 2.30 8.34 2.58 ;
        RECT  8.12 2.30 8.28 3.48 ;
        RECT  7.02 2.30 7.30 2.58 ;
        RECT  7.08 2.30 7.24 3.48 ;
        RECT  6.14 2.52 6.42 3.48 ;
        RECT  4.06 2.52 4.34 3.48 ;
        RECT  1.74 1.92 2.02 2.20 ;
        RECT  1.80 1.92 1.96 3.48 ;
        RECT  0.62 1.84 0.90 2.12 ;
        RECT  0.68 1.84 0.84 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 8.80 0.28 ;
        RECT  8.12 -0.28 8.62 0.32 ;
        RECT  8.06 0.58 8.34 0.86 ;
        RECT  8.12 -0.28 8.28 0.86 ;
        RECT  7.02 0.58 7.30 0.86 ;
        RECT  7.08 -0.28 7.24 0.86 ;
        RECT  5.90 0.72 6.18 1.00 ;
        RECT  5.96 -0.28 6.12 1.00 ;
        RECT  3.82 0.72 4.10 1.00 ;
        RECT  3.88 -0.28 4.04 1.00 ;
        RECT  1.74 0.72 2.02 1.00 ;
        RECT  1.80 -0.28 1.96 1.00 ;
        RECT  0.62 0.52 0.90 0.80 ;
        RECT  0.68 -0.28 0.84 0.80 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.08 0.52 0.38 0.80 ;
        RECT  0.08 1.01 1.10 1.17 ;
        RECT  0.82 0.96 1.10 1.24 ;
        RECT  0.08 0.52 0.24 2.12 ;
        RECT  0.08 1.84 0.38 2.12 ;
        RECT  1.14 0.52 1.42 0.80 ;
        RECT  1.26 1.40 1.56 1.68 ;
        RECT  1.26 0.52 1.42 2.12 ;
        RECT  1.14 1.84 1.42 2.12 ;
        RECT  2.26 0.72 2.54 1.00 ;
        RECT  2.32 0.72 2.48 2.20 ;
        RECT  2.26 1.92 2.54 2.20 ;
        RECT  3.24 0.72 3.58 1.00 ;
        RECT  3.24 0.72 3.40 2.20 ;
        RECT  3.24 1.92 3.58 2.20 ;
        RECT  2.78 0.72 3.06 1.00 ;
        RECT  4.04 1.48 4.32 1.76 ;
        RECT  3.74 1.60 4.32 1.76 ;
        RECT  2.84 0.72 3.00 2.20 ;
        RECT  2.78 1.92 3.06 2.20 ;
        RECT  2.90 1.92 3.06 2.52 ;
        RECT  3.74 1.60 3.90 2.52 ;
        RECT  2.90 2.36 3.90 2.52 ;
        RECT  4.34 0.72 4.64 1.00 ;
        RECT  3.56 1.16 4.64 1.32 ;
        RECT  3.56 1.16 3.84 1.44 ;
        RECT  4.48 0.72 4.64 2.20 ;
        RECT  4.34 1.92 4.64 2.20 ;
        RECT  5.32 0.72 5.66 1.00 ;
        RECT  5.32 0.72 5.48 2.20 ;
        RECT  5.32 1.92 5.66 2.20 ;
        RECT  4.86 0.72 5.14 1.00 ;
        RECT  6.12 1.48 6.40 1.76 ;
        RECT  5.82 1.60 6.40 1.76 ;
        RECT  4.92 0.72 5.08 2.20 ;
        RECT  4.86 1.92 5.14 2.20 ;
        RECT  4.98 1.92 5.14 2.52 ;
        RECT  5.82 1.60 5.98 2.52 ;
        RECT  4.98 2.36 5.98 2.52 ;
        RECT  6.42 0.72 6.72 1.00 ;
        RECT  5.64 1.16 6.72 1.32 ;
        RECT  5.64 1.16 5.92 1.44 ;
        RECT  6.56 1.54 7.48 1.70 ;
        RECT  7.20 1.48 7.48 1.76 ;
        RECT  6.56 0.72 6.72 2.20 ;
        RECT  6.42 1.92 6.72 2.20 ;
    END
END DFFSSP4V1_0

MACRO DFFSSP2V1_1
    CLASS CORE ;
    FOREIGN DFFSSP2V1_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 14.89  LAYER ME1  ;
        ANTENNADIFFAREA 6.69  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.55  LAYER ME1  ;
        ANTENNAMAXAREACAR 27.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.66 1.46 7.92 1.74 ;
        RECT  7.60 1.84 7.88 2.12 ;
        RECT  7.66 0.96 7.88 2.12 ;
        RECT  7.60 0.96 7.88 1.24 ;
        END
    END Q
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.88 1.39 1.16 1.81 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.39 0.72 1.81 ;
        END
    END D
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 8.00 0.28 ;
        RECT  7.54 -0.28 7.82 0.32 ;
        RECT  7.08 0.64 7.36 0.92 ;
        RECT  7.14 -0.28 7.30 0.92 ;
        RECT  6.08 0.96 6.36 1.24 ;
        RECT  6.18 -0.28 6.34 1.24 ;
        RECT  3.36 0.72 3.64 1.00 ;
        RECT  3.42 -0.28 3.58 1.00 ;
        RECT  0.62 0.68 0.90 0.96 ;
        RECT  0.68 -0.28 0.84 0.96 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 8.00 3.48 ;
        RECT  7.54 2.88 7.82 3.48 ;
        RECT  7.08 2.16 7.36 2.44 ;
        RECT  7.14 2.16 7.30 3.48 ;
        RECT  6.08 2.62 6.36 3.48 ;
        RECT  3.48 1.92 3.76 2.20 ;
        RECT  3.54 1.92 3.70 3.48 ;
        RECT  0.38 2.62 0.66 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  1.14 0.68 1.48 0.96 ;
        RECT  1.32 1.22 1.64 1.50 ;
        RECT  1.32 0.68 1.48 2.25 ;
        RECT  1.14 1.97 1.48 2.25 ;
        RECT  0.08 0.68 0.38 0.96 ;
        RECT  1.68 0.72 1.96 1.00 ;
        RECT  0.08 0.68 0.24 2.25 ;
        RECT  0.08 1.97 0.38 2.25 ;
        RECT  1.80 0.72 1.96 2.20 ;
        RECT  0.08 2.09 0.98 2.25 ;
        RECT  0.82 2.09 0.98 2.57 ;
        RECT  1.68 1.92 1.84 2.57 ;
        RECT  0.82 2.41 1.84 2.57 ;
        RECT  2.76 0.72 3.07 1.00 ;
        RECT  2.76 0.72 2.92 2.20 ;
        RECT  2.72 1.92 3.00 2.20 ;
        RECT  2.20 0.72 2.48 1.00 ;
        RECT  3.56 1.48 3.84 1.76 ;
        RECT  3.16 1.60 3.84 1.76 ;
        RECT  2.26 0.72 2.42 2.20 ;
        RECT  2.20 1.92 2.48 2.20 ;
        RECT  2.32 1.92 2.48 2.52 ;
        RECT  3.16 1.60 3.32 2.52 ;
        RECT  2.32 2.36 3.32 2.52 ;
        RECT  3.88 0.72 4.16 1.00 ;
        RECT  3.08 1.16 4.16 1.32 ;
        RECT  3.08 1.16 3.36 1.44 ;
        RECT  4.00 0.72 4.16 2.20 ;
        RECT  4.00 1.92 4.28 2.20 ;
        RECT  4.56 0.44 6.02 0.60 ;
        RECT  5.74 0.44 6.02 0.80 ;
        RECT  4.44 0.76 4.72 1.04 ;
        RECT  4.56 0.44 4.72 2.20 ;
        RECT  4.52 1.92 4.80 2.20 ;
        RECT  5.56 0.96 5.84 1.24 ;
        RECT  5.56 1.46 6.56 1.62 ;
        RECT  6.28 1.40 6.56 1.68 ;
        RECT  5.56 0.96 5.72 2.12 ;
        RECT  5.56 1.84 5.84 2.12 ;
        RECT  4.96 0.76 5.24 1.04 ;
        RECT  6.60 0.96 6.88 1.24 ;
        RECT  6.60 1.84 6.88 2.12 ;
        RECT  5.08 0.76 5.24 2.20 ;
        RECT  5.04 1.92 5.32 2.20 ;
        RECT  5.16 1.92 5.32 2.44 ;
        RECT  6.72 0.96 6.88 2.44 ;
        RECT  5.16 2.28 6.88 2.44 ;
    END
END DFFSSP2V1_1

MACRO DFFSSP2V1_0
    CLASS CORE ;
    FOREIGN DFFSSP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 14.86  LAYER ME1  ;
        ANTENNADIFFAREA 7.05  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.79  LAYER ME1  ;
        ANTENNAMAXAREACAR 18.88  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.54 1.92 7.88 2.20 ;
        RECT  7.72 0.96 7.88 2.20 ;
        RECT  7.54 0.96 7.88 1.24 ;
        END
    END Q
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.40 0.82 1.68 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.72 1.40 2.14 1.68 ;
        END
    END D
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 8.00 0.28 ;
        RECT  7.54 -0.28 7.82 0.32 ;
        RECT  7.02 0.62 7.30 0.90 ;
        RECT  7.08 -0.28 7.24 0.90 ;
        RECT  5.90 0.72 6.18 1.00 ;
        RECT  5.96 -0.28 6.12 1.00 ;
        RECT  3.82 0.72 4.10 1.00 ;
        RECT  3.88 -0.28 4.04 1.00 ;
        RECT  1.74 0.72 2.02 1.00 ;
        RECT  1.80 -0.28 1.96 1.00 ;
        RECT  0.62 0.52 0.90 0.80 ;
        RECT  0.68 -0.28 0.84 0.80 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 8.00 3.48 ;
        RECT  7.54 2.88 7.82 3.48 ;
        RECT  7.02 2.26 7.30 2.54 ;
        RECT  7.08 2.26 7.24 3.48 ;
        RECT  6.14 2.52 6.42 3.48 ;
        RECT  4.06 2.52 4.34 3.48 ;
        RECT  1.74 1.92 2.02 2.20 ;
        RECT  1.80 1.92 1.96 3.48 ;
        RECT  0.62 1.84 0.90 2.12 ;
        RECT  0.68 1.84 0.84 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.08 0.52 0.38 0.80 ;
        RECT  0.08 1.01 1.10 1.17 ;
        RECT  0.82 0.96 1.10 1.24 ;
        RECT  0.08 0.52 0.24 2.12 ;
        RECT  0.08 1.84 0.38 2.12 ;
        RECT  1.14 0.52 1.42 0.80 ;
        RECT  1.26 1.40 1.56 1.68 ;
        RECT  1.26 0.52 1.42 2.12 ;
        RECT  1.14 1.84 1.42 2.12 ;
        RECT  2.26 0.72 2.54 1.00 ;
        RECT  2.32 0.72 2.48 2.20 ;
        RECT  2.26 1.92 2.54 2.20 ;
        RECT  3.24 0.72 3.58 1.00 ;
        RECT  3.24 0.72 3.40 2.20 ;
        RECT  3.24 1.92 3.58 2.20 ;
        RECT  2.78 0.72 3.06 1.00 ;
        RECT  4.04 1.48 4.32 1.76 ;
        RECT  3.74 1.60 4.32 1.76 ;
        RECT  2.84 0.72 3.00 2.20 ;
        RECT  2.78 1.92 3.06 2.20 ;
        RECT  2.90 1.92 3.06 2.52 ;
        RECT  3.74 1.60 3.90 2.52 ;
        RECT  2.90 2.36 3.90 2.52 ;
        RECT  4.34 0.72 4.64 1.00 ;
        RECT  3.56 1.16 4.64 1.32 ;
        RECT  3.56 1.16 3.84 1.44 ;
        RECT  4.48 0.72 4.64 2.20 ;
        RECT  4.34 1.92 4.64 2.20 ;
        RECT  5.32 0.72 5.66 1.00 ;
        RECT  5.32 0.72 5.48 2.20 ;
        RECT  5.32 1.92 5.66 2.20 ;
        RECT  4.86 0.72 5.14 1.00 ;
        RECT  6.12 1.48 6.40 1.76 ;
        RECT  5.82 1.60 6.40 1.76 ;
        RECT  4.92 0.72 5.08 2.20 ;
        RECT  4.86 1.92 5.14 2.20 ;
        RECT  4.98 1.92 5.14 2.52 ;
        RECT  5.82 1.60 5.98 2.52 ;
        RECT  4.98 2.36 5.98 2.52 ;
        RECT  6.42 0.72 6.72 1.00 ;
        RECT  5.64 1.16 6.72 1.32 ;
        RECT  5.64 1.16 5.92 1.44 ;
        RECT  6.56 1.54 7.48 1.70 ;
        RECT  7.20 1.48 7.48 1.76 ;
        RECT  6.56 0.72 6.72 2.20 ;
        RECT  6.42 1.92 6.72 2.20 ;
    END
END DFFSSP2V1_0

MACRO DFFSSP1V1_1
    CLASS CORE ;
    FOREIGN DFFSSP1V1_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.39 0.72 1.81 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.88 1.39 1.16 1.81 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 14.99  LAYER ME1  ;
        ANTENNADIFFAREA 6.25  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.47  LAYER ME1  ;
        ANTENNAMAXAREACAR 31.86  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.66 1.46 7.92 1.74 ;
        RECT  7.60 1.84 7.88 2.12 ;
        RECT  7.66 0.96 7.88 2.12 ;
        RECT  7.60 0.96 7.88 1.24 ;
        END
    END Q
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 8.00 3.48 ;
        RECT  7.54 2.88 7.82 3.48 ;
        RECT  7.08 1.84 7.36 2.12 ;
        RECT  7.14 1.84 7.30 3.48 ;
        RECT  6.08 2.62 6.36 3.48 ;
        RECT  3.48 1.92 3.76 2.20 ;
        RECT  3.54 1.92 3.70 3.48 ;
        RECT  0.38 2.62 0.66 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 8.00 0.28 ;
        RECT  7.54 -0.28 7.82 0.32 ;
        RECT  7.08 0.96 7.36 1.24 ;
        RECT  7.14 -0.28 7.30 1.24 ;
        RECT  6.08 0.96 6.36 1.24 ;
        RECT  6.18 -0.28 6.34 1.24 ;
        RECT  3.36 0.72 3.64 1.00 ;
        RECT  3.42 -0.28 3.58 1.00 ;
        RECT  0.62 0.68 0.90 0.96 ;
        RECT  0.68 -0.28 0.84 0.96 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  1.14 0.68 1.48 0.96 ;
        RECT  1.32 1.22 1.64 1.50 ;
        RECT  1.32 0.68 1.48 2.25 ;
        RECT  1.14 1.97 1.48 2.25 ;
        RECT  0.08 0.68 0.38 0.96 ;
        RECT  1.68 0.72 1.96 1.00 ;
        RECT  0.08 0.68 0.24 2.25 ;
        RECT  0.08 1.97 0.38 2.25 ;
        RECT  1.80 0.72 1.96 2.20 ;
        RECT  0.08 2.09 0.98 2.25 ;
        RECT  0.82 2.09 0.98 2.57 ;
        RECT  1.68 1.92 1.84 2.57 ;
        RECT  0.82 2.41 1.84 2.57 ;
        RECT  2.76 0.72 3.07 1.00 ;
        RECT  2.76 0.72 2.92 2.20 ;
        RECT  2.72 1.92 3.00 2.20 ;
        RECT  2.20 0.72 2.48 1.00 ;
        RECT  3.56 1.48 3.84 1.76 ;
        RECT  3.16 1.60 3.84 1.76 ;
        RECT  2.26 0.72 2.42 2.20 ;
        RECT  2.20 1.92 2.48 2.20 ;
        RECT  2.32 1.92 2.48 2.52 ;
        RECT  3.16 1.60 3.32 2.52 ;
        RECT  2.32 2.36 3.32 2.52 ;
        RECT  3.88 0.72 4.16 1.00 ;
        RECT  3.08 1.16 4.16 1.32 ;
        RECT  3.08 1.16 3.36 1.44 ;
        RECT  4.00 0.72 4.16 2.20 ;
        RECT  4.00 1.92 4.28 2.20 ;
        RECT  4.56 0.44 6.02 0.60 ;
        RECT  5.74 0.44 6.02 0.80 ;
        RECT  4.44 0.76 4.72 1.04 ;
        RECT  4.56 0.44 4.72 2.20 ;
        RECT  4.52 1.92 4.80 2.20 ;
        RECT  5.56 0.96 5.84 1.24 ;
        RECT  5.56 1.46 6.56 1.62 ;
        RECT  6.28 1.40 6.56 1.68 ;
        RECT  5.56 0.96 5.72 2.12 ;
        RECT  5.56 1.84 5.84 2.12 ;
        RECT  4.96 0.76 5.24 1.04 ;
        RECT  6.60 0.96 6.88 1.24 ;
        RECT  6.60 1.84 6.88 2.12 ;
        RECT  5.08 0.76 5.24 2.20 ;
        RECT  5.04 1.92 5.32 2.20 ;
        RECT  5.16 1.92 5.32 2.44 ;
        RECT  6.72 0.96 6.88 2.44 ;
        RECT  5.16 2.28 6.88 2.44 ;
    END
END DFFSSP1V1_1

MACRO DFFSSP1V1_0
    CLASS CORE ;
    FOREIGN DFFSSP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.72 1.40 2.14 1.68 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.40 0.82 1.68 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 14.97  LAYER ME1  ;
        ANTENNADIFFAREA 6.59  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.71  LAYER ME1  ;
        ANTENNAMAXAREACAR 21.21  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.54 1.92 7.88 2.20 ;
        RECT  7.72 0.96 7.88 2.20 ;
        RECT  7.54 0.96 7.88 1.24 ;
        END
    END Q
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 8.00 3.48 ;
        RECT  7.54 2.88 7.82 3.48 ;
        RECT  7.02 1.92 7.30 2.20 ;
        RECT  7.08 1.92 7.24 3.48 ;
        RECT  6.14 2.52 6.42 3.48 ;
        RECT  4.06 2.52 4.34 3.48 ;
        RECT  1.74 1.92 2.02 2.20 ;
        RECT  1.80 1.92 1.96 3.48 ;
        RECT  0.62 1.84 0.90 2.12 ;
        RECT  0.68 1.84 0.84 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 8.00 0.28 ;
        RECT  7.54 -0.28 7.82 0.32 ;
        RECT  7.02 0.96 7.30 1.24 ;
        RECT  7.08 -0.28 7.24 1.24 ;
        RECT  5.90 0.72 6.18 1.00 ;
        RECT  5.96 -0.28 6.12 1.00 ;
        RECT  3.82 0.72 4.10 1.00 ;
        RECT  3.88 -0.28 4.04 1.00 ;
        RECT  1.74 0.72 2.02 1.00 ;
        RECT  1.80 -0.28 1.96 1.00 ;
        RECT  0.62 0.52 0.90 0.80 ;
        RECT  0.68 -0.28 0.84 0.80 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.08 0.52 0.38 0.80 ;
        RECT  0.08 1.01 1.10 1.17 ;
        RECT  0.82 0.96 1.10 1.24 ;
        RECT  0.08 0.52 0.24 2.12 ;
        RECT  0.08 1.84 0.38 2.12 ;
        RECT  1.14 0.52 1.42 0.80 ;
        RECT  1.26 1.40 1.56 1.68 ;
        RECT  1.26 0.52 1.42 2.12 ;
        RECT  1.14 1.84 1.42 2.12 ;
        RECT  2.26 0.72 2.54 1.00 ;
        RECT  2.32 0.72 2.48 2.20 ;
        RECT  2.26 1.92 2.54 2.20 ;
        RECT  3.24 0.72 3.58 1.00 ;
        RECT  3.24 0.72 3.40 2.20 ;
        RECT  3.24 1.92 3.58 2.20 ;
        RECT  2.78 0.72 3.06 1.00 ;
        RECT  4.04 1.48 4.32 1.76 ;
        RECT  3.74 1.60 4.32 1.76 ;
        RECT  2.84 0.72 3.00 2.20 ;
        RECT  2.78 1.92 3.06 2.20 ;
        RECT  2.90 1.92 3.06 2.52 ;
        RECT  3.74 1.60 3.90 2.52 ;
        RECT  2.90 2.36 3.90 2.52 ;
        RECT  4.34 0.72 4.64 1.00 ;
        RECT  3.56 1.16 4.64 1.32 ;
        RECT  3.56 1.16 3.84 1.44 ;
        RECT  4.48 0.72 4.64 2.20 ;
        RECT  4.34 1.92 4.64 2.20 ;
        RECT  5.32 0.72 5.66 1.00 ;
        RECT  5.32 0.72 5.48 2.20 ;
        RECT  5.32 1.92 5.66 2.20 ;
        RECT  4.86 0.72 5.14 1.00 ;
        RECT  6.12 1.48 6.40 1.76 ;
        RECT  5.82 1.60 6.40 1.76 ;
        RECT  4.92 0.72 5.08 2.20 ;
        RECT  4.86 1.92 5.14 2.20 ;
        RECT  4.98 1.92 5.14 2.52 ;
        RECT  5.82 1.60 5.98 2.52 ;
        RECT  4.98 2.36 5.98 2.52 ;
        RECT  6.42 0.72 6.72 1.00 ;
        RECT  5.64 1.16 6.72 1.32 ;
        RECT  5.64 1.16 5.92 1.44 ;
        RECT  6.56 1.54 7.48 1.70 ;
        RECT  7.20 1.48 7.48 1.76 ;
        RECT  6.56 0.72 6.72 2.20 ;
        RECT  6.42 1.92 6.72 2.20 ;
    END
END DFFSSP1V1_0

MACRO DFFSRZSP8V1_0
    CLASS CORE ;
    FOREIGN DFFSRZSP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 26.12  LAYER ME1  ;
        ANTENNADIFFAREA 12.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.05  LAYER ME1  ;
        ANTENNAMAXAREACAR 24.96  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.83 1.90 13.11 2.50 ;
        RECT  12.83 0.64 13.11 1.24 ;
        RECT  12.83 0.64 12.99 2.50 ;
        RECT  11.66 1.52 12.99 1.68 ;
        RECT  11.79 1.90 12.07 2.50 ;
        RECT  11.79 0.64 12.07 1.24 ;
        RECT  11.79 0.64 11.95 2.50 ;
        RECT  11.66 1.46 11.95 1.74 ;
        END
    END Q
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.21 1.40 3.53 1.76 ;
        END
    END CK
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.22 1.40 9.60 1.68 ;
        END
    END RB
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.87  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 12.90  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.06 1.46 2.34 1.74 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.81 2.23 2.25 ;
        RECT  1.95 0.81 2.23 1.09 ;
        END
    END TD
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END SEL
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.20  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.83  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.81 1.19 2.25 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  0.91 0.81 1.19 1.09 ;
        END
    END D
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 14.00 0.28 ;
        RECT  13.41 -0.28 13.82 0.32 ;
        RECT  13.35 0.64 13.63 1.24 ;
        RECT  13.41 -0.28 13.57 1.24 ;
        RECT  12.31 0.64 12.59 1.24 ;
        RECT  12.37 -0.28 12.53 1.24 ;
        RECT  11.27 0.64 11.55 1.24 ;
        RECT  11.33 -0.28 11.49 1.24 ;
        RECT  10.27 0.88 10.55 1.16 ;
        RECT  10.33 -0.28 10.49 1.16 ;
        RECT  7.29 -0.28 7.57 0.72 ;
        RECT  2.71 -0.28 2.99 0.68 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 14.00 3.48 ;
        RECT  13.41 2.88 13.82 3.48 ;
        RECT  13.35 1.90 13.63 2.50 ;
        RECT  13.41 1.90 13.57 3.48 ;
        RECT  12.31 1.90 12.59 2.50 ;
        RECT  12.37 1.90 12.53 3.48 ;
        RECT  11.27 1.90 11.55 2.50 ;
        RECT  11.33 1.90 11.49 3.48 ;
        RECT  10.27 1.84 10.55 2.12 ;
        RECT  10.33 1.84 10.49 3.48 ;
        RECT  9.23 1.84 9.51 2.12 ;
        RECT  9.29 1.84 9.45 3.48 ;
        RECT  8.39 1.84 8.55 3.48 ;
        RECT  8.19 1.84 8.55 2.12 ;
        RECT  2.71 2.52 2.99 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  1.55 1.97 1.71 2.57 ;
        RECT  1.55 2.41 2.37 2.57 ;
        RECT  2.09 2.41 2.37 2.69 ;
        RECT  3.47 0.96 3.85 1.24 ;
        RECT  3.69 1.46 3.97 1.74 ;
        RECT  3.69 0.96 3.85 2.20 ;
        RECT  3.47 1.92 3.85 2.20 ;
        RECT  4.07 0.44 4.35 0.72 ;
        RECT  3.15 0.56 4.35 0.72 ;
        RECT  3.15 0.56 3.31 1.12 ;
        RECT  2.43 0.96 3.31 1.12 ;
        RECT  2.43 0.96 2.71 1.24 ;
        RECT  2.50 0.96 2.66 2.20 ;
        RECT  2.43 1.92 2.71 2.20 ;
        RECT  2.43 2.04 3.31 2.20 ;
        RECT  3.15 2.04 3.31 2.64 ;
        RECT  3.15 2.48 4.35 2.64 ;
        RECT  4.07 2.48 4.35 2.76 ;
        RECT  5.67 0.88 5.95 1.16 ;
        RECT  5.67 0.88 5.83 2.12 ;
        RECT  5.45 1.84 5.83 2.12 ;
        RECT  6.15 1.84 6.43 2.12 ;
        RECT  5.45 1.96 6.43 2.12 ;
        RECT  6.85 0.44 7.13 0.72 ;
        RECT  6.31 0.56 7.13 0.72 ;
        RECT  6.19 0.88 6.47 1.16 ;
        RECT  6.31 0.56 6.47 1.68 ;
        RECT  6.31 1.52 6.75 1.68 ;
        RECT  6.59 1.52 6.75 2.12 ;
        RECT  6.59 1.84 6.95 2.12 ;
        RECT  4.63 0.87 4.91 1.15 ;
        RECT  4.07 0.99 4.91 1.15 ;
        RECT  4.07 0.96 4.35 1.24 ;
        RECT  4.19 0.96 4.35 2.12 ;
        RECT  4.19 1.84 4.47 2.12 ;
        RECT  4.19 1.96 4.77 2.12 ;
        RECT  4.61 1.96 4.77 2.76 ;
        RECT  7.95 2.42 8.23 2.76 ;
        RECT  4.61 2.60 8.23 2.76 ;
        RECT  8.15 0.50 8.43 0.78 ;
        RECT  6.71 0.88 6.99 1.20 ;
        RECT  7.33 0.92 7.61 1.20 ;
        RECT  8.15 0.50 8.31 1.20 ;
        RECT  6.71 1.04 8.31 1.20 ;
        RECT  7.11 1.04 7.27 2.12 ;
        RECT  7.11 1.84 7.47 2.12 ;
        RECT  5.13 0.87 5.43 1.15 ;
        RECT  8.81 0.92 9.09 1.20 ;
        RECT  7.63 1.52 8.97 1.68 ;
        RECT  8.81 0.92 8.97 2.12 ;
        RECT  5.01 1.84 5.29 2.12 ;
        RECT  8.71 1.84 8.99 2.12 ;
        RECT  5.13 0.87 5.29 2.44 ;
        RECT  7.63 1.52 7.79 2.44 ;
        RECT  5.13 2.28 7.79 2.44 ;
        RECT  9.37 0.88 9.65 1.16 ;
        RECT  9.37 1.00 9.92 1.16 ;
        RECT  9.76 1.46 10.75 1.62 ;
        RECT  10.47 1.40 10.75 1.68 ;
        RECT  9.76 1.00 9.92 2.12 ;
        RECT  9.75 1.84 10.03 2.12 ;
        RECT  10.79 0.88 11.07 1.16 ;
        RECT  10.79 1.84 11.07 2.12 ;
        RECT  10.91 0.88 11.07 2.76 ;
        RECT  10.82 2.48 11.10 2.76 ;
    END
END DFFSRZSP8V1_0

MACRO DFFSRZSP4V1_0
    CLASS CORE ;
    FOREIGN DFFSRZSP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.20  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.83  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.81 1.19 2.25 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  0.91 0.81 1.19 1.09 ;
        END
    END D
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END SEL
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.87  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 12.90  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.06 1.46 2.34 1.74 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.81 2.23 2.25 ;
        RECT  1.95 0.81 2.23 1.09 ;
        END
    END TD
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.22 1.40 9.60 1.68 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.21 1.40 3.53 1.76 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 23.72  LAYER ME1  ;
        ANTENNADIFFAREA 10.17  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.76  LAYER ME1  ;
        ANTENNAMAXAREACAR 31.28  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.79 1.90 12.07 2.50 ;
        RECT  11.79 0.64 12.07 1.24 ;
        RECT  11.79 0.64 11.95 2.50 ;
        RECT  11.66 1.46 11.95 1.74 ;
        END
    END Q
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 12.80 3.48 ;
        RECT  12.34 2.88 12.62 3.48 ;
        RECT  12.31 1.90 12.59 2.50 ;
        RECT  12.37 1.90 12.53 3.48 ;
        RECT  11.27 1.90 11.55 2.50 ;
        RECT  11.33 1.90 11.49 3.48 ;
        RECT  10.27 1.84 10.55 2.12 ;
        RECT  10.33 1.84 10.49 3.48 ;
        RECT  9.23 1.84 9.51 2.12 ;
        RECT  9.29 1.84 9.45 3.48 ;
        RECT  8.39 1.84 8.55 3.48 ;
        RECT  8.19 1.84 8.55 2.12 ;
        RECT  2.71 2.52 2.99 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 12.80 0.28 ;
        RECT  12.34 -0.28 12.62 0.32 ;
        RECT  12.31 0.64 12.59 1.24 ;
        RECT  12.37 -0.28 12.53 1.24 ;
        RECT  11.27 0.64 11.55 1.24 ;
        RECT  11.33 -0.28 11.49 1.24 ;
        RECT  10.27 0.88 10.55 1.16 ;
        RECT  10.33 -0.28 10.49 1.16 ;
        RECT  7.29 -0.28 7.57 0.72 ;
        RECT  2.71 -0.28 2.99 0.68 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  1.55 1.97 1.71 2.57 ;
        RECT  1.55 2.41 2.37 2.57 ;
        RECT  2.09 2.41 2.37 2.69 ;
        RECT  3.47 0.96 3.85 1.24 ;
        RECT  3.69 1.46 3.97 1.74 ;
        RECT  3.69 0.96 3.85 2.20 ;
        RECT  3.47 1.92 3.85 2.20 ;
        RECT  4.07 0.44 4.35 0.72 ;
        RECT  3.15 0.56 4.35 0.72 ;
        RECT  3.15 0.56 3.31 1.12 ;
        RECT  2.43 0.96 3.31 1.12 ;
        RECT  2.43 0.96 2.71 1.24 ;
        RECT  2.50 0.96 2.66 2.20 ;
        RECT  2.43 1.92 2.71 2.20 ;
        RECT  2.43 2.04 3.31 2.20 ;
        RECT  3.15 2.04 3.31 2.64 ;
        RECT  3.15 2.48 4.35 2.64 ;
        RECT  4.07 2.48 4.35 2.76 ;
        RECT  5.67 0.88 5.95 1.16 ;
        RECT  5.67 0.88 5.83 2.12 ;
        RECT  5.45 1.84 5.83 2.12 ;
        RECT  6.15 1.84 6.43 2.12 ;
        RECT  5.45 1.96 6.43 2.12 ;
        RECT  6.85 0.44 7.13 0.72 ;
        RECT  6.31 0.56 7.13 0.72 ;
        RECT  6.19 0.88 6.47 1.16 ;
        RECT  6.31 0.56 6.47 1.68 ;
        RECT  6.31 1.52 6.75 1.68 ;
        RECT  6.59 1.52 6.75 2.12 ;
        RECT  6.59 1.84 6.95 2.12 ;
        RECT  4.63 0.87 4.91 1.15 ;
        RECT  4.07 0.99 4.91 1.15 ;
        RECT  4.07 0.96 4.35 1.24 ;
        RECT  4.19 0.96 4.35 2.12 ;
        RECT  4.19 1.84 4.47 2.12 ;
        RECT  4.19 1.96 4.77 2.12 ;
        RECT  4.61 1.96 4.77 2.76 ;
        RECT  7.95 2.42 8.23 2.76 ;
        RECT  4.61 2.60 8.23 2.76 ;
        RECT  8.15 0.50 8.43 0.78 ;
        RECT  6.71 0.88 6.99 1.20 ;
        RECT  7.33 0.92 7.61 1.20 ;
        RECT  8.15 0.50 8.31 1.20 ;
        RECT  6.71 1.04 8.31 1.20 ;
        RECT  7.11 1.04 7.27 2.12 ;
        RECT  7.11 1.84 7.47 2.12 ;
        RECT  5.13 0.87 5.43 1.15 ;
        RECT  8.81 0.92 9.09 1.20 ;
        RECT  7.63 1.52 8.97 1.68 ;
        RECT  8.81 0.92 8.97 2.12 ;
        RECT  5.01 1.84 5.29 2.12 ;
        RECT  8.71 1.84 8.99 2.12 ;
        RECT  5.13 0.87 5.29 2.44 ;
        RECT  7.63 1.52 7.79 2.44 ;
        RECT  5.13 2.28 7.79 2.44 ;
        RECT  9.37 0.88 9.65 1.16 ;
        RECT  9.37 1.00 9.92 1.16 ;
        RECT  9.76 1.46 10.75 1.62 ;
        RECT  10.47 1.40 10.75 1.68 ;
        RECT  9.76 1.00 9.92 2.12 ;
        RECT  9.75 1.84 10.03 2.12 ;
        RECT  10.79 0.88 11.07 1.16 ;
        RECT  10.79 1.84 11.07 2.12 ;
        RECT  10.91 0.88 11.07 2.76 ;
        RECT  10.82 2.48 11.10 2.76 ;
    END
END DFFSRZSP4V1_0

MACRO DFFSRZSP2V1_0
    CLASS CORE ;
    FOREIGN DFFSRZSP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 22.82  LAYER ME1  ;
        ANTENNADIFFAREA 9.57  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.61  LAYER ME1  ;
        ANTENNAMAXAREACAR 37.15  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.79 1.90 12.07 2.50 ;
        RECT  11.79 0.64 12.07 1.24 ;
        RECT  11.79 0.64 11.95 2.50 ;
        RECT  11.66 1.46 11.95 1.74 ;
        END
    END Q
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.21 1.40 3.53 1.76 ;
        END
    END CK
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.22 1.40 9.60 1.68 ;
        END
    END RB
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.87  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 12.90  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.06 1.46 2.34 1.74 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.81 2.23 2.25 ;
        RECT  1.95 0.81 2.23 1.09 ;
        END
    END TD
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END SEL
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.20  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.83  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.81 1.19 2.25 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  0.91 0.81 1.19 1.09 ;
        END
    END D
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 12.40 0.28 ;
        RECT  11.94 -0.28 12.22 0.32 ;
        RECT  11.27 0.64 11.55 1.24 ;
        RECT  11.33 -0.28 11.49 1.24 ;
        RECT  10.27 0.88 10.55 1.16 ;
        RECT  10.33 -0.28 10.49 1.16 ;
        RECT  7.29 -0.28 7.57 0.72 ;
        RECT  2.71 -0.28 2.99 0.68 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 12.40 3.48 ;
        RECT  11.94 2.88 12.22 3.48 ;
        RECT  11.27 1.90 11.55 2.50 ;
        RECT  11.33 1.90 11.49 3.48 ;
        RECT  10.27 1.84 10.55 2.12 ;
        RECT  10.33 1.84 10.49 3.48 ;
        RECT  9.23 1.84 9.51 2.12 ;
        RECT  9.29 1.84 9.45 3.48 ;
        RECT  8.39 1.84 8.55 3.48 ;
        RECT  8.19 1.84 8.55 2.12 ;
        RECT  2.71 2.52 2.99 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  1.55 1.97 1.71 2.57 ;
        RECT  1.55 2.41 2.37 2.57 ;
        RECT  2.09 2.41 2.37 2.69 ;
        RECT  3.47 0.96 3.85 1.24 ;
        RECT  3.69 1.46 3.97 1.74 ;
        RECT  3.69 0.96 3.85 2.20 ;
        RECT  3.47 1.92 3.85 2.20 ;
        RECT  4.07 0.44 4.35 0.72 ;
        RECT  3.15 0.56 4.35 0.72 ;
        RECT  3.15 0.56 3.31 1.12 ;
        RECT  2.43 0.96 3.31 1.12 ;
        RECT  2.43 0.96 2.71 1.24 ;
        RECT  2.50 0.96 2.66 2.20 ;
        RECT  2.43 1.92 2.71 2.20 ;
        RECT  2.43 2.04 3.31 2.20 ;
        RECT  3.15 2.04 3.31 2.64 ;
        RECT  3.15 2.48 4.35 2.64 ;
        RECT  4.07 2.48 4.35 2.76 ;
        RECT  5.67 0.88 5.95 1.16 ;
        RECT  5.67 0.88 5.83 2.12 ;
        RECT  5.45 1.84 5.83 2.12 ;
        RECT  6.15 1.84 6.43 2.12 ;
        RECT  5.45 1.96 6.43 2.12 ;
        RECT  6.85 0.44 7.13 0.72 ;
        RECT  6.31 0.56 7.13 0.72 ;
        RECT  6.19 0.88 6.47 1.16 ;
        RECT  6.31 0.56 6.47 1.68 ;
        RECT  6.31 1.52 6.75 1.68 ;
        RECT  6.59 1.52 6.75 2.12 ;
        RECT  6.59 1.84 6.95 2.12 ;
        RECT  4.63 0.87 4.91 1.15 ;
        RECT  4.07 0.99 4.91 1.15 ;
        RECT  4.07 0.96 4.35 1.24 ;
        RECT  4.19 0.96 4.35 2.12 ;
        RECT  4.19 1.84 4.47 2.12 ;
        RECT  4.19 1.96 4.77 2.12 ;
        RECT  4.61 1.96 4.77 2.76 ;
        RECT  7.95 2.42 8.23 2.76 ;
        RECT  4.61 2.60 8.23 2.76 ;
        RECT  8.15 0.50 8.43 0.78 ;
        RECT  6.71 0.88 6.99 1.20 ;
        RECT  7.33 0.92 7.61 1.20 ;
        RECT  8.15 0.50 8.31 1.20 ;
        RECT  6.71 1.04 8.31 1.20 ;
        RECT  7.11 1.04 7.27 2.12 ;
        RECT  7.11 1.84 7.47 2.12 ;
        RECT  5.13 0.87 5.43 1.15 ;
        RECT  8.81 0.92 9.09 1.20 ;
        RECT  7.63 1.52 8.97 1.68 ;
        RECT  8.81 0.92 8.97 2.12 ;
        RECT  5.01 1.84 5.29 2.12 ;
        RECT  8.71 1.84 8.99 2.12 ;
        RECT  5.13 0.87 5.29 2.44 ;
        RECT  7.63 1.52 7.79 2.44 ;
        RECT  5.13 2.28 7.79 2.44 ;
        RECT  9.37 0.88 9.65 1.16 ;
        RECT  9.37 1.00 9.92 1.16 ;
        RECT  9.76 1.46 10.75 1.62 ;
        RECT  10.47 1.40 10.75 1.68 ;
        RECT  9.76 1.00 9.92 2.12 ;
        RECT  9.75 1.84 10.03 2.12 ;
        RECT  10.79 0.88 11.07 1.16 ;
        RECT  10.79 1.84 11.07 2.12 ;
        RECT  10.91 0.88 11.07 2.76 ;
        RECT  10.82 2.48 11.10 2.76 ;
    END
END DFFSRZSP2V1_0

MACRO DFFSRZSP1V1_0
    CLASS CORE ;
    FOREIGN DFFSRZSP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.20  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.83  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.81 1.19 2.25 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  0.91 0.81 1.19 1.09 ;
        END
    END D
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END SEL
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.87  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 12.90  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.06 1.46 2.34 1.74 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.81 2.23 2.25 ;
        RECT  1.95 0.81 2.23 1.09 ;
        END
    END TD
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.22 1.40 9.60 1.68 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.21 1.40 3.53 1.76 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 22.26  LAYER ME1  ;
        ANTENNADIFFAREA 9.13  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.54  LAYER ME1  ;
        ANTENNAMAXAREACAR 41.40  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.79 1.90 12.07 2.18 ;
        RECT  11.79 0.88 12.07 1.16 ;
        RECT  11.79 0.88 11.95 2.18 ;
        RECT  11.66 1.46 11.95 1.74 ;
        END
    END Q
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 12.40 3.48 ;
        RECT  11.94 2.88 12.22 3.48 ;
        RECT  11.27 1.90 11.55 2.18 ;
        RECT  11.33 1.90 11.49 3.48 ;
        RECT  10.27 1.84 10.55 2.12 ;
        RECT  10.33 1.84 10.49 3.48 ;
        RECT  9.23 1.84 9.51 2.12 ;
        RECT  9.29 1.84 9.45 3.48 ;
        RECT  8.39 1.84 8.55 3.48 ;
        RECT  8.19 1.84 8.55 2.12 ;
        RECT  2.71 2.52 2.99 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 12.40 0.28 ;
        RECT  11.94 -0.28 12.22 0.32 ;
        RECT  11.27 0.88 11.55 1.16 ;
        RECT  11.33 -0.28 11.49 1.16 ;
        RECT  10.27 0.88 10.55 1.16 ;
        RECT  10.33 -0.28 10.49 1.16 ;
        RECT  7.29 -0.28 7.57 0.72 ;
        RECT  2.71 -0.28 2.99 0.68 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  1.55 1.97 1.71 2.57 ;
        RECT  1.55 2.41 2.37 2.57 ;
        RECT  2.09 2.41 2.37 2.69 ;
        RECT  3.47 0.96 3.85 1.24 ;
        RECT  3.69 1.46 3.97 1.74 ;
        RECT  3.69 0.96 3.85 2.20 ;
        RECT  3.47 1.92 3.85 2.20 ;
        RECT  4.07 0.44 4.35 0.72 ;
        RECT  3.15 0.56 4.35 0.72 ;
        RECT  3.15 0.56 3.31 1.12 ;
        RECT  2.43 0.96 3.31 1.12 ;
        RECT  2.43 0.96 2.71 1.24 ;
        RECT  2.50 0.96 2.66 2.20 ;
        RECT  2.43 1.92 2.71 2.20 ;
        RECT  2.43 2.04 3.31 2.20 ;
        RECT  3.15 2.04 3.31 2.64 ;
        RECT  3.15 2.48 4.35 2.64 ;
        RECT  4.07 2.48 4.35 2.76 ;
        RECT  5.67 0.88 5.95 1.16 ;
        RECT  5.67 0.88 5.83 2.12 ;
        RECT  5.45 1.84 5.83 2.12 ;
        RECT  6.15 1.84 6.43 2.12 ;
        RECT  5.45 1.96 6.43 2.12 ;
        RECT  6.85 0.44 7.13 0.72 ;
        RECT  6.31 0.56 7.13 0.72 ;
        RECT  6.19 0.88 6.47 1.16 ;
        RECT  6.31 0.56 6.47 1.68 ;
        RECT  6.31 1.52 6.75 1.68 ;
        RECT  6.59 1.52 6.75 2.12 ;
        RECT  6.59 1.84 6.95 2.12 ;
        RECT  4.63 0.87 4.91 1.15 ;
        RECT  4.07 0.99 4.91 1.15 ;
        RECT  4.07 0.96 4.35 1.24 ;
        RECT  4.19 0.96 4.35 2.12 ;
        RECT  4.19 1.84 4.47 2.12 ;
        RECT  4.19 1.96 4.77 2.12 ;
        RECT  4.61 1.96 4.77 2.76 ;
        RECT  7.95 2.42 8.23 2.76 ;
        RECT  4.61 2.60 8.23 2.76 ;
        RECT  8.15 0.50 8.43 0.78 ;
        RECT  6.71 0.88 6.99 1.20 ;
        RECT  7.33 0.92 7.61 1.20 ;
        RECT  8.15 0.50 8.31 1.20 ;
        RECT  6.71 1.04 8.31 1.20 ;
        RECT  7.11 1.04 7.27 2.12 ;
        RECT  7.11 1.84 7.47 2.12 ;
        RECT  5.13 0.87 5.43 1.15 ;
        RECT  8.81 0.92 9.09 1.20 ;
        RECT  7.63 1.52 8.97 1.68 ;
        RECT  8.81 0.92 8.97 2.12 ;
        RECT  5.01 1.84 5.29 2.12 ;
        RECT  8.71 1.84 8.99 2.12 ;
        RECT  5.13 0.87 5.29 2.44 ;
        RECT  7.63 1.52 7.79 2.44 ;
        RECT  5.13 2.28 7.79 2.44 ;
        RECT  9.37 0.88 9.65 1.16 ;
        RECT  9.37 1.00 9.92 1.16 ;
        RECT  9.76 1.46 10.75 1.62 ;
        RECT  10.47 1.40 10.75 1.68 ;
        RECT  9.76 1.00 9.92 2.12 ;
        RECT  9.75 1.84 10.03 2.12 ;
        RECT  10.79 0.88 11.07 1.16 ;
        RECT  10.79 1.84 11.07 2.12 ;
        RECT  10.91 0.88 11.07 2.76 ;
        RECT  10.82 2.48 11.10 2.76 ;
    END
END DFFSRZSP1V1_0

MACRO DFFSRSZSP8V1_0
    CLASS CORE ;
    FOREIGN DFFSRSZSP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 28.77  LAYER ME1  ;
        ANTENNADIFFAREA 13.38  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.05  LAYER ME1  ;
        ANTENNAMAXAREACAR 27.49  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.47 1.90 14.75 2.50 ;
        RECT  14.47 0.64 14.75 1.24 ;
        RECT  14.47 0.64 14.63 2.50 ;
        RECT  13.55 1.52 14.63 1.68 ;
        RECT  13.55 1.46 13.94 1.74 ;
        RECT  13.43 1.90 13.71 2.50 ;
        RECT  13.55 0.64 13.71 2.50 ;
        RECT  13.43 0.64 13.71 1.24 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.66 0.44 11.94 0.94 ;
        RECT  11.45 0.44 11.94 0.72 ;
        END
    END SB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.99 1.40 10.41 1.68 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.24 1.40 3.54 1.76 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.87  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 12.90  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.06 1.46 2.34 1.74 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.81 2.23 2.25 ;
        RECT  1.95 0.81 2.23 1.09 ;
        END
    END TD
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END SEL
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.20  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.83  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.81 1.19 2.25 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  0.91 0.81 1.19 1.09 ;
        END
    END D
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 15.60 0.28 ;
        RECT  15.05 -0.28 15.42 0.32 ;
        RECT  14.99 0.64 15.27 1.24 ;
        RECT  15.05 -0.28 15.21 1.24 ;
        RECT  13.95 0.64 14.23 1.24 ;
        RECT  14.01 -0.28 14.17 1.24 ;
        RECT  12.91 0.64 13.19 1.24 ;
        RECT  12.97 -0.28 13.13 1.24 ;
        RECT  11.08 0.88 11.43 1.16 ;
        RECT  11.08 -0.28 11.24 1.16 ;
        RECT  8.69 -0.28 8.97 0.68 ;
        RECT  2.71 -0.28 2.99 0.68 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 15.60 3.48 ;
        RECT  15.05 2.88 15.42 3.48 ;
        RECT  14.99 1.90 15.27 2.50 ;
        RECT  15.05 1.90 15.21 3.48 ;
        RECT  13.95 1.90 14.23 2.50 ;
        RECT  14.01 1.90 14.17 3.48 ;
        RECT  12.91 1.90 13.19 2.50 ;
        RECT  12.97 1.90 13.13 3.48 ;
        RECT  12.31 2.40 12.59 3.48 ;
        RECT  11.09 1.84 11.37 2.12 ;
        RECT  11.15 1.84 11.31 3.48 ;
        RECT  10.05 1.84 10.33 2.12 ;
        RECT  10.11 1.84 10.27 3.48 ;
        RECT  8.77 1.96 9.29 2.12 ;
        RECT  9.01 1.84 9.29 2.12 ;
        RECT  8.65 2.52 8.93 3.48 ;
        RECT  8.77 1.96 8.93 3.48 ;
        RECT  2.71 2.52 2.99 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  1.55 1.97 1.71 2.57 ;
        RECT  1.55 2.41 2.37 2.57 ;
        RECT  2.09 2.41 2.37 2.69 ;
        RECT  3.47 0.96 3.86 1.24 ;
        RECT  3.70 1.46 4.02 1.74 ;
        RECT  3.70 0.96 3.86 2.20 ;
        RECT  3.47 1.92 3.86 2.20 ;
        RECT  4.07 0.44 4.35 0.72 ;
        RECT  3.15 0.56 4.35 0.72 ;
        RECT  3.15 0.56 3.31 1.12 ;
        RECT  2.43 0.96 3.31 1.12 ;
        RECT  2.43 0.96 2.71 1.24 ;
        RECT  2.55 0.96 2.71 2.20 ;
        RECT  2.43 1.92 2.71 2.20 ;
        RECT  2.43 2.04 3.31 2.20 ;
        RECT  3.15 2.04 3.31 2.64 ;
        RECT  3.15 2.48 4.25 2.64 ;
        RECT  3.97 2.48 4.25 2.76 ;
        RECT  5.59 0.88 5.91 1.16 ;
        RECT  5.59 0.88 5.75 2.00 ;
        RECT  5.25 1.84 6.23 2.00 ;
        RECT  5.25 1.84 5.53 2.12 ;
        RECT  5.95 1.84 6.23 2.12 ;
        RECT  6.15 0.88 6.43 1.16 ;
        RECT  6.27 0.88 6.43 1.58 ;
        RECT  7.11 1.14 7.39 1.58 ;
        RECT  6.27 1.42 7.39 1.58 ;
        RECT  6.39 1.42 6.55 2.12 ;
        RECT  6.39 1.84 6.75 2.12 ;
        RECT  4.75 0.50 8.15 0.66 ;
        RECT  7.87 0.50 8.15 0.78 ;
        RECT  4.63 0.86 4.91 1.14 ;
        RECT  4.75 0.50 4.91 1.14 ;
        RECT  4.07 0.98 4.91 1.14 ;
        RECT  4.07 0.96 4.35 1.24 ;
        RECT  4.29 0.98 4.45 2.12 ;
        RECT  4.29 1.84 4.57 2.12 ;
        RECT  9.13 0.50 9.41 0.78 ;
        RECT  6.67 0.82 7.71 0.98 ;
        RECT  6.67 0.82 6.95 1.16 ;
        RECT  9.13 0.50 9.29 1.16 ;
        RECT  7.55 1.00 9.29 1.16 ;
        RECT  7.55 0.96 7.91 1.24 ;
        RECT  7.85 1.00 8.01 2.12 ;
        RECT  6.99 1.84 7.27 2.12 ;
        RECT  7.85 1.84 8.19 2.12 ;
        RECT  6.99 1.96 8.19 2.12 ;
        RECT  5.07 0.86 5.43 1.14 ;
        RECT  9.67 0.96 10.11 1.24 ;
        RECT  5.07 0.86 5.23 1.48 ;
        RECT  8.35 1.52 9.83 1.68 ;
        RECT  4.81 1.84 5.09 2.12 ;
        RECT  9.67 0.96 9.83 2.12 ;
        RECT  9.53 1.84 9.83 2.12 ;
        RECT  4.93 1.32 5.09 2.44 ;
        RECT  8.35 1.52 8.51 2.44 ;
        RECT  4.93 2.28 8.51 2.44 ;
        RECT  10.31 0.88 10.73 1.16 ;
        RECT  10.57 1.46 12.11 1.62 ;
        RECT  11.83 1.40 12.11 1.68 ;
        RECT  10.57 0.88 10.73 2.12 ;
        RECT  10.57 1.84 10.85 2.12 ;
        RECT  12.11 0.88 12.47 1.16 ;
        RECT  12.31 0.88 12.47 2.16 ;
        RECT  11.82 1.96 12.59 2.12 ;
        RECT  12.31 1.88 12.59 2.16 ;
        RECT  11.82 1.96 11.98 2.76 ;
        RECT  11.70 2.48 11.98 2.76 ;
    END
END DFFSRSZSP8V1_0

MACRO DFFSRSZSP4V1_0
    CLASS CORE ;
    FOREIGN DFFSRSZSP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.20  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.83  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.81 1.19 2.25 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  0.91 0.81 1.19 1.09 ;
        END
    END D
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END SEL
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.87  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 12.90  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.06 1.46 2.34 1.74 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.81 2.23 2.25 ;
        RECT  1.95 0.81 2.23 1.09 ;
        END
    END TD
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.24 1.40 3.54 1.76 ;
        END
    END CK
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.99 1.40 10.41 1.68 ;
        END
    END RB
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.66 0.44 11.94 0.94 ;
        RECT  11.45 0.44 11.94 0.72 ;
        END
    END SB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 26.43  LAYER ME1  ;
        ANTENNADIFFAREA 11.56  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.76  LAYER ME1  ;
        ANTENNAMAXAREACAR 34.85  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.55 1.46 13.94 1.74 ;
        RECT  13.43 1.90 13.71 2.50 ;
        RECT  13.55 0.64 13.71 2.50 ;
        RECT  13.43 0.64 13.71 1.24 ;
        END
    END Q
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 14.40 3.48 ;
        RECT  13.95 1.90 14.23 2.50 ;
        RECT  13.94 2.88 14.22 3.48 ;
        RECT  14.01 1.90 14.17 3.48 ;
        RECT  12.91 1.90 13.19 2.50 ;
        RECT  12.97 1.90 13.13 3.48 ;
        RECT  12.31 2.40 12.59 3.48 ;
        RECT  11.09 1.84 11.37 2.12 ;
        RECT  11.15 1.84 11.31 3.48 ;
        RECT  10.05 1.84 10.33 2.12 ;
        RECT  10.11 1.84 10.27 3.48 ;
        RECT  8.77 1.96 9.29 2.12 ;
        RECT  9.01 1.84 9.29 2.12 ;
        RECT  8.65 2.52 8.93 3.48 ;
        RECT  8.77 1.96 8.93 3.48 ;
        RECT  2.71 2.52 2.99 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 14.40 0.28 ;
        RECT  13.95 0.64 14.23 1.24 ;
        RECT  13.94 -0.28 14.22 0.32 ;
        RECT  14.01 -0.28 14.17 1.24 ;
        RECT  12.91 0.64 13.19 1.24 ;
        RECT  12.97 -0.28 13.13 1.24 ;
        RECT  11.08 0.88 11.43 1.16 ;
        RECT  11.08 -0.28 11.24 1.16 ;
        RECT  8.69 -0.28 8.97 0.68 ;
        RECT  2.71 -0.28 2.99 0.68 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  1.55 1.97 1.71 2.57 ;
        RECT  1.55 2.41 2.37 2.57 ;
        RECT  2.09 2.41 2.37 2.69 ;
        RECT  3.47 0.96 3.86 1.24 ;
        RECT  3.70 1.46 4.02 1.74 ;
        RECT  3.70 0.96 3.86 2.20 ;
        RECT  3.47 1.92 3.86 2.20 ;
        RECT  4.07 0.44 4.35 0.72 ;
        RECT  3.15 0.56 4.35 0.72 ;
        RECT  3.15 0.56 3.31 1.12 ;
        RECT  2.43 0.96 3.31 1.12 ;
        RECT  2.43 0.96 2.71 1.24 ;
        RECT  2.55 0.96 2.71 2.20 ;
        RECT  2.43 1.92 2.71 2.20 ;
        RECT  2.43 2.04 3.31 2.20 ;
        RECT  3.15 2.04 3.31 2.64 ;
        RECT  3.15 2.48 4.25 2.64 ;
        RECT  3.97 2.48 4.25 2.76 ;
        RECT  5.59 0.88 5.91 1.16 ;
        RECT  5.59 0.88 5.75 2.00 ;
        RECT  5.25 1.84 6.23 2.00 ;
        RECT  5.25 1.84 5.53 2.12 ;
        RECT  5.95 1.84 6.23 2.12 ;
        RECT  6.15 0.88 6.43 1.16 ;
        RECT  6.27 0.88 6.43 1.58 ;
        RECT  7.11 1.14 7.39 1.58 ;
        RECT  6.27 1.42 7.39 1.58 ;
        RECT  6.39 1.42 6.55 2.12 ;
        RECT  6.39 1.84 6.75 2.12 ;
        RECT  4.75 0.50 8.15 0.66 ;
        RECT  7.87 0.50 8.15 0.78 ;
        RECT  4.63 0.86 4.91 1.14 ;
        RECT  4.75 0.50 4.91 1.14 ;
        RECT  4.07 0.98 4.91 1.14 ;
        RECT  4.07 0.96 4.35 1.24 ;
        RECT  4.29 0.98 4.45 2.12 ;
        RECT  4.29 1.84 4.57 2.12 ;
        RECT  9.13 0.50 9.41 0.78 ;
        RECT  6.67 0.82 7.71 0.98 ;
        RECT  6.67 0.82 6.95 1.16 ;
        RECT  9.13 0.50 9.29 1.16 ;
        RECT  7.55 1.00 9.29 1.16 ;
        RECT  7.55 0.96 7.91 1.24 ;
        RECT  7.85 1.00 8.01 2.12 ;
        RECT  6.99 1.84 7.27 2.12 ;
        RECT  7.85 1.84 8.19 2.12 ;
        RECT  6.99 1.96 8.19 2.12 ;
        RECT  5.07 0.86 5.43 1.14 ;
        RECT  9.67 0.96 10.11 1.24 ;
        RECT  5.07 0.86 5.23 1.48 ;
        RECT  8.35 1.52 9.83 1.68 ;
        RECT  4.81 1.84 5.09 2.12 ;
        RECT  9.67 0.96 9.83 2.12 ;
        RECT  9.53 1.84 9.83 2.12 ;
        RECT  4.93 1.32 5.09 2.44 ;
        RECT  8.35 1.52 8.51 2.44 ;
        RECT  4.93 2.28 8.51 2.44 ;
        RECT  10.31 0.88 10.73 1.16 ;
        RECT  10.57 1.46 12.11 1.62 ;
        RECT  11.83 1.40 12.11 1.68 ;
        RECT  10.57 0.88 10.73 2.12 ;
        RECT  10.57 1.84 10.85 2.12 ;
        RECT  12.11 0.88 12.47 1.16 ;
        RECT  12.31 0.88 12.47 2.16 ;
        RECT  11.82 1.96 12.59 2.12 ;
        RECT  12.31 1.88 12.59 2.16 ;
        RECT  11.82 1.96 11.98 2.76 ;
        RECT  11.70 2.48 11.98 2.76 ;
    END
END DFFSRSZSP4V1_0

MACRO DFFSRSZSP2V1_0
    CLASS CORE ;
    FOREIGN DFFSRSZSP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 25.53  LAYER ME1  ;
        ANTENNADIFFAREA 10.95  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.61  LAYER ME1  ;
        ANTENNAMAXAREACAR 41.55  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.55 1.46 13.92 1.74 ;
        RECT  13.43 1.90 13.71 2.50 ;
        RECT  13.55 0.64 13.71 2.50 ;
        RECT  13.43 0.64 13.71 1.24 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.66 0.44 11.94 0.94 ;
        RECT  11.45 0.44 11.94 0.72 ;
        END
    END SB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.99 1.40 10.41 1.68 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.24 1.40 3.54 1.76 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.87  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 12.90  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.06 1.46 2.34 1.74 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.81 2.23 2.25 ;
        RECT  1.95 0.81 2.23 1.09 ;
        END
    END TD
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END SEL
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.20  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.83  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.81 1.19 2.25 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  0.91 0.81 1.19 1.09 ;
        END
    END D
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 14.00 0.28 ;
        RECT  13.54 -0.28 13.82 0.32 ;
        RECT  12.91 0.64 13.19 1.24 ;
        RECT  12.97 -0.28 13.13 1.24 ;
        RECT  11.08 0.88 11.43 1.16 ;
        RECT  11.08 -0.28 11.24 1.16 ;
        RECT  8.69 -0.28 8.97 0.68 ;
        RECT  2.71 -0.28 2.99 0.68 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 14.00 3.48 ;
        RECT  13.54 2.88 13.82 3.48 ;
        RECT  12.91 1.90 13.19 2.50 ;
        RECT  12.97 1.90 13.13 3.48 ;
        RECT  12.31 2.40 12.59 3.48 ;
        RECT  11.09 1.84 11.37 2.12 ;
        RECT  11.15 1.84 11.31 3.48 ;
        RECT  10.05 1.84 10.33 2.12 ;
        RECT  10.11 1.84 10.27 3.48 ;
        RECT  8.77 1.96 9.29 2.12 ;
        RECT  9.01 1.84 9.29 2.12 ;
        RECT  8.65 2.52 8.93 3.48 ;
        RECT  8.77 1.96 8.93 3.48 ;
        RECT  2.71 2.52 2.99 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  1.55 1.97 1.71 2.57 ;
        RECT  1.55 2.41 2.37 2.57 ;
        RECT  2.09 2.41 2.37 2.69 ;
        RECT  3.47 0.96 3.86 1.24 ;
        RECT  3.70 1.46 4.02 1.74 ;
        RECT  3.70 0.96 3.86 2.20 ;
        RECT  3.47 1.92 3.86 2.20 ;
        RECT  4.07 0.44 4.35 0.72 ;
        RECT  3.15 0.56 4.35 0.72 ;
        RECT  3.15 0.56 3.31 1.12 ;
        RECT  2.43 0.96 3.31 1.12 ;
        RECT  2.43 0.96 2.71 1.24 ;
        RECT  2.55 0.96 2.71 2.20 ;
        RECT  2.43 1.92 2.71 2.20 ;
        RECT  2.43 2.04 3.31 2.20 ;
        RECT  3.15 2.04 3.31 2.64 ;
        RECT  3.15 2.48 4.25 2.64 ;
        RECT  3.97 2.48 4.25 2.76 ;
        RECT  5.59 0.88 5.91 1.16 ;
        RECT  5.59 0.88 5.75 2.00 ;
        RECT  5.25 1.84 6.23 2.00 ;
        RECT  5.25 1.84 5.53 2.12 ;
        RECT  5.95 1.84 6.23 2.12 ;
        RECT  6.15 0.88 6.43 1.16 ;
        RECT  6.27 0.88 6.43 1.58 ;
        RECT  7.11 1.14 7.39 1.58 ;
        RECT  6.27 1.42 7.39 1.58 ;
        RECT  6.39 1.42 6.55 2.12 ;
        RECT  6.39 1.84 6.75 2.12 ;
        RECT  4.75 0.50 8.15 0.66 ;
        RECT  7.87 0.50 8.15 0.78 ;
        RECT  4.63 0.86 4.91 1.14 ;
        RECT  4.75 0.50 4.91 1.14 ;
        RECT  4.07 0.98 4.91 1.14 ;
        RECT  4.07 0.96 4.35 1.24 ;
        RECT  4.29 0.98 4.45 2.12 ;
        RECT  4.29 1.84 4.57 2.12 ;
        RECT  9.13 0.50 9.41 0.78 ;
        RECT  6.67 0.82 7.71 0.98 ;
        RECT  6.67 0.82 6.95 1.16 ;
        RECT  9.13 0.50 9.29 1.16 ;
        RECT  7.55 1.00 9.29 1.16 ;
        RECT  7.55 0.96 7.91 1.24 ;
        RECT  7.85 1.00 8.01 2.12 ;
        RECT  6.99 1.84 7.27 2.12 ;
        RECT  7.85 1.84 8.19 2.12 ;
        RECT  6.99 1.96 8.19 2.12 ;
        RECT  5.07 0.86 5.43 1.14 ;
        RECT  9.67 0.96 10.11 1.24 ;
        RECT  5.07 0.86 5.23 1.48 ;
        RECT  8.35 1.52 9.83 1.68 ;
        RECT  4.81 1.84 5.09 2.12 ;
        RECT  9.67 0.96 9.83 2.12 ;
        RECT  9.53 1.84 9.83 2.12 ;
        RECT  4.93 1.32 5.09 2.44 ;
        RECT  8.35 1.52 8.51 2.44 ;
        RECT  4.93 2.28 8.51 2.44 ;
        RECT  10.31 0.88 10.73 1.16 ;
        RECT  10.57 1.46 12.11 1.62 ;
        RECT  11.83 1.40 12.11 1.68 ;
        RECT  10.57 0.88 10.73 2.12 ;
        RECT  10.57 1.84 10.85 2.12 ;
        RECT  12.11 0.88 12.47 1.16 ;
        RECT  12.31 0.88 12.47 2.16 ;
        RECT  11.82 1.96 12.59 2.12 ;
        RECT  12.31 1.88 12.59 2.16 ;
        RECT  11.82 1.96 11.98 2.76 ;
        RECT  11.70 2.48 11.98 2.76 ;
    END
END DFFSRSZSP2V1_0

MACRO DFFSRSZSP1V1_0
    CLASS CORE ;
    FOREIGN DFFSRSZSP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.66 0.44 11.94 0.94 ;
        RECT  11.45 0.44 11.94 0.72 ;
        END
    END SB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.99 1.40 10.41 1.68 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.24 1.40 3.54 1.76 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 24.95  LAYER ME1  ;
        ANTENNADIFFAREA 10.52  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.54  LAYER ME1  ;
        ANTENNAMAXAREACAR 46.41  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.55 1.46 13.92 1.74 ;
        RECT  13.43 1.90 13.71 2.18 ;
        RECT  13.55 0.96 13.71 2.18 ;
        RECT  13.43 0.96 13.71 1.24 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.20  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.83  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.81 1.19 2.25 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  0.91 0.81 1.19 1.09 ;
        END
    END D
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.87  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 12.90  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.06 1.46 2.34 1.74 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.81 2.23 2.25 ;
        RECT  1.95 0.81 2.23 1.09 ;
        END
    END TD
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END SEL
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 14.00 3.48 ;
        RECT  13.54 2.88 13.82 3.48 ;
        RECT  12.91 1.90 13.19 2.18 ;
        RECT  12.97 1.90 13.13 3.48 ;
        RECT  12.31 2.40 12.59 3.48 ;
        RECT  11.09 1.84 11.37 2.12 ;
        RECT  11.15 1.84 11.31 3.48 ;
        RECT  10.05 1.84 10.33 2.12 ;
        RECT  10.11 1.84 10.27 3.48 ;
        RECT  8.77 1.96 9.29 2.12 ;
        RECT  9.01 1.84 9.29 2.12 ;
        RECT  8.65 2.52 8.93 3.48 ;
        RECT  8.77 1.96 8.93 3.48 ;
        RECT  2.71 2.52 2.99 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 14.00 0.28 ;
        RECT  13.54 -0.28 13.82 0.32 ;
        RECT  12.91 0.96 13.19 1.24 ;
        RECT  12.97 -0.28 13.13 1.24 ;
        RECT  11.08 0.88 11.43 1.16 ;
        RECT  11.08 -0.28 11.24 1.16 ;
        RECT  8.69 -0.28 8.97 0.68 ;
        RECT  2.71 -0.28 2.99 0.68 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  1.55 1.97 1.71 2.57 ;
        RECT  1.55 2.41 2.37 2.57 ;
        RECT  2.09 2.41 2.37 2.69 ;
        RECT  3.47 0.96 3.86 1.24 ;
        RECT  3.70 1.46 4.02 1.74 ;
        RECT  3.70 0.96 3.86 2.20 ;
        RECT  3.47 1.92 3.86 2.20 ;
        RECT  4.07 0.44 4.35 0.72 ;
        RECT  3.15 0.56 4.35 0.72 ;
        RECT  3.15 0.56 3.31 1.12 ;
        RECT  2.43 0.96 3.31 1.12 ;
        RECT  2.43 0.96 2.71 1.24 ;
        RECT  2.55 0.96 2.71 2.20 ;
        RECT  2.43 1.92 2.71 2.20 ;
        RECT  2.43 2.04 3.31 2.20 ;
        RECT  3.15 2.04 3.31 2.64 ;
        RECT  3.15 2.48 4.25 2.64 ;
        RECT  3.97 2.48 4.25 2.76 ;
        RECT  5.59 0.88 5.91 1.16 ;
        RECT  5.59 0.88 5.75 2.00 ;
        RECT  5.25 1.84 6.23 2.00 ;
        RECT  5.25 1.84 5.53 2.12 ;
        RECT  5.95 1.84 6.23 2.12 ;
        RECT  6.15 0.88 6.43 1.16 ;
        RECT  6.27 0.88 6.43 1.58 ;
        RECT  7.11 1.14 7.39 1.58 ;
        RECT  6.27 1.42 7.39 1.58 ;
        RECT  6.39 1.42 6.55 2.12 ;
        RECT  6.39 1.84 6.75 2.12 ;
        RECT  4.75 0.50 8.15 0.66 ;
        RECT  7.87 0.50 8.15 0.78 ;
        RECT  4.63 0.86 4.91 1.14 ;
        RECT  4.75 0.50 4.91 1.14 ;
        RECT  4.07 0.98 4.91 1.14 ;
        RECT  4.07 0.96 4.35 1.24 ;
        RECT  4.29 0.98 4.45 2.12 ;
        RECT  4.29 1.84 4.57 2.12 ;
        RECT  9.13 0.50 9.41 0.78 ;
        RECT  6.67 0.82 7.71 0.98 ;
        RECT  6.67 0.82 6.95 1.16 ;
        RECT  9.13 0.50 9.29 1.16 ;
        RECT  7.55 1.00 9.29 1.16 ;
        RECT  7.55 0.96 7.91 1.24 ;
        RECT  7.85 1.00 8.01 2.12 ;
        RECT  6.99 1.84 7.27 2.12 ;
        RECT  7.85 1.84 8.19 2.12 ;
        RECT  6.99 1.96 8.19 2.12 ;
        RECT  5.07 0.86 5.43 1.14 ;
        RECT  9.67 0.96 10.11 1.24 ;
        RECT  5.07 0.86 5.23 1.48 ;
        RECT  8.35 1.52 9.83 1.68 ;
        RECT  4.81 1.84 5.09 2.12 ;
        RECT  9.67 0.96 9.83 2.12 ;
        RECT  9.53 1.84 9.83 2.12 ;
        RECT  4.93 1.32 5.09 2.44 ;
        RECT  8.35 1.52 8.51 2.44 ;
        RECT  4.93 2.28 8.51 2.44 ;
        RECT  10.31 0.88 10.73 1.16 ;
        RECT  10.57 1.46 12.11 1.62 ;
        RECT  11.83 1.40 12.11 1.68 ;
        RECT  10.57 0.88 10.73 2.12 ;
        RECT  10.57 1.84 10.85 2.12 ;
        RECT  12.11 0.88 12.47 1.16 ;
        RECT  12.31 0.88 12.47 2.16 ;
        RECT  11.82 1.96 12.59 2.12 ;
        RECT  12.31 1.88 12.59 2.16 ;
        RECT  11.82 1.96 11.98 2.76 ;
        RECT  11.70 2.48 11.98 2.76 ;
    END
END DFFSRSZSP1V1_0

MACRO DFFSRSSP8V1_0
    CLASS CORE ;
    FOREIGN DFFSRSSP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 13.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 25.48  LAYER ME1  ;
        ANTENNADIFFAREA 12.23  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.98  LAYER ME1  ;
        ANTENNAMAXAREACAR 26.02  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.14 1.88 12.42 2.48 ;
        RECT  12.14 0.64 12.42 1.24 ;
        RECT  12.14 0.64 12.30 2.48 ;
        RECT  11.22 1.52 12.30 1.68 ;
        RECT  11.22 1.46 11.54 1.74 ;
        RECT  11.10 1.88 11.38 2.48 ;
        RECT  11.22 0.64 11.38 2.48 ;
        RECT  11.10 0.64 11.38 1.24 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.40 0.70 1.76 ;
        END
    END D
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.66 1.40 8.08 1.68 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.40 1.16 1.76 ;
        END
    END CK
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.26 0.44 9.54 0.94 ;
        RECT  9.07 0.44 9.54 0.72 ;
        END
    END SB
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 13.20 3.48 ;
        RECT  12.72 2.88 13.02 3.48 ;
        RECT  12.66 1.88 12.94 2.48 ;
        RECT  12.72 1.88 12.88 3.48 ;
        RECT  11.62 1.88 11.90 2.48 ;
        RECT  11.68 1.88 11.84 3.48 ;
        RECT  10.58 1.88 10.86 2.48 ;
        RECT  10.64 1.88 10.80 3.48 ;
        RECT  9.98 2.40 10.26 3.48 ;
        RECT  8.76 1.84 9.04 2.12 ;
        RECT  8.82 1.84 8.98 3.48 ;
        RECT  7.72 1.84 8.00 2.12 ;
        RECT  7.78 1.84 7.94 3.48 ;
        RECT  6.44 1.96 6.96 2.12 ;
        RECT  6.68 1.84 6.96 2.12 ;
        RECT  6.32 2.52 6.60 3.48 ;
        RECT  6.44 1.96 6.60 3.48 ;
        RECT  0.38 2.48 0.66 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 13.20 0.28 ;
        RECT  12.72 -0.28 13.02 0.32 ;
        RECT  12.66 0.64 12.94 1.24 ;
        RECT  12.72 -0.28 12.88 1.24 ;
        RECT  11.62 0.64 11.90 1.24 ;
        RECT  11.68 -0.28 11.84 1.24 ;
        RECT  10.58 0.64 10.86 1.24 ;
        RECT  10.64 -0.28 10.80 1.24 ;
        RECT  8.75 0.88 9.10 1.16 ;
        RECT  8.75 -0.28 8.91 1.16 ;
        RECT  6.36 -0.28 6.64 0.68 ;
        RECT  0.38 -0.28 0.66 0.68 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  1.14 0.96 1.48 1.24 ;
        RECT  1.32 1.46 1.64 1.74 ;
        RECT  1.32 0.96 1.48 2.20 ;
        RECT  1.14 1.92 1.48 2.20 ;
        RECT  1.74 0.44 2.02 0.72 ;
        RECT  0.82 0.56 2.02 0.72 ;
        RECT  0.82 0.56 0.98 1.12 ;
        RECT  0.08 0.96 0.98 1.12 ;
        RECT  0.08 0.96 0.38 1.24 ;
        RECT  0.08 0.96 0.24 2.20 ;
        RECT  0.08 1.92 0.38 2.20 ;
        RECT  0.08 2.04 0.98 2.20 ;
        RECT  0.82 2.04 0.98 2.64 ;
        RECT  0.82 2.48 1.92 2.64 ;
        RECT  1.64 2.48 1.92 2.76 ;
        RECT  3.26 0.88 3.58 1.16 ;
        RECT  3.26 0.88 3.42 2.00 ;
        RECT  2.92 1.84 3.90 2.00 ;
        RECT  2.92 1.84 3.20 2.12 ;
        RECT  3.62 1.84 3.90 2.12 ;
        RECT  3.82 0.88 4.10 1.16 ;
        RECT  3.94 0.88 4.10 1.58 ;
        RECT  4.78 1.14 5.06 1.58 ;
        RECT  3.94 1.42 5.06 1.58 ;
        RECT  4.06 1.42 4.22 2.12 ;
        RECT  4.06 1.84 4.42 2.12 ;
        RECT  2.42 0.50 5.82 0.66 ;
        RECT  5.54 0.50 5.82 0.78 ;
        RECT  2.30 0.86 2.58 1.14 ;
        RECT  2.42 0.50 2.58 1.14 ;
        RECT  1.74 0.98 2.58 1.14 ;
        RECT  1.74 0.96 2.02 1.24 ;
        RECT  1.96 0.98 2.12 2.12 ;
        RECT  1.96 1.84 2.24 2.12 ;
        RECT  6.80 0.50 7.08 0.78 ;
        RECT  4.34 0.82 5.38 0.98 ;
        RECT  4.34 0.82 4.62 1.16 ;
        RECT  6.80 0.50 6.96 1.16 ;
        RECT  5.22 1.00 6.96 1.16 ;
        RECT  5.22 0.96 5.58 1.24 ;
        RECT  5.52 1.00 5.68 2.12 ;
        RECT  4.66 1.84 4.94 2.12 ;
        RECT  5.52 1.84 5.86 2.12 ;
        RECT  4.66 1.96 5.86 2.12 ;
        RECT  2.74 0.86 3.10 1.14 ;
        RECT  7.34 0.96 7.78 1.24 ;
        RECT  2.74 0.86 2.90 1.48 ;
        RECT  6.02 1.52 7.50 1.68 ;
        RECT  2.48 1.84 2.76 2.12 ;
        RECT  7.34 0.96 7.50 2.12 ;
        RECT  7.20 1.84 7.50 2.12 ;
        RECT  2.60 1.32 2.76 2.44 ;
        RECT  6.02 1.52 6.18 2.44 ;
        RECT  2.60 2.28 6.18 2.44 ;
        RECT  7.98 0.88 8.40 1.16 ;
        RECT  8.24 1.46 9.78 1.62 ;
        RECT  9.50 1.40 9.78 1.68 ;
        RECT  8.24 0.88 8.40 2.12 ;
        RECT  8.24 1.84 8.52 2.12 ;
        RECT  9.78 0.88 10.14 1.16 ;
        RECT  9.98 0.88 10.14 2.16 ;
        RECT  9.49 1.96 10.26 2.12 ;
        RECT  9.98 1.88 10.26 2.16 ;
        RECT  9.49 1.96 9.65 2.76 ;
        RECT  9.37 2.48 9.65 2.76 ;
    END
END DFFSRSSP8V1_0

MACRO DFFSRSSP4V1_0
    CLASS CORE ;
    FOREIGN DFFSRSSP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.26 0.44 9.54 0.94 ;
        RECT  9.07 0.44 9.54 0.72 ;
        END
    END SB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.40 1.16 1.76 ;
        END
    END CK
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.66 1.40 8.08 1.68 ;
        END
    END RB
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.40 0.70 1.76 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 23.13  LAYER ME1  ;
        ANTENNADIFFAREA 10.40  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.69  LAYER ME1  ;
        ANTENNAMAXAREACAR 33.46  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.22 1.46 11.54 1.74 ;
        RECT  11.10 1.90 11.38 2.50 ;
        RECT  11.22 0.64 11.38 2.50 ;
        RECT  11.10 0.64 11.38 1.24 ;
        END
    END Q
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 12.00 3.48 ;
        RECT  11.62 1.90 11.90 2.50 ;
        RECT  11.54 2.88 11.84 3.48 ;
        RECT  11.68 1.90 11.84 3.48 ;
        RECT  10.58 1.90 10.86 2.50 ;
        RECT  10.64 1.90 10.80 3.48 ;
        RECT  9.98 2.40 10.26 3.48 ;
        RECT  8.76 1.84 9.04 2.12 ;
        RECT  8.82 1.84 8.98 3.48 ;
        RECT  7.72 1.84 8.00 2.12 ;
        RECT  7.78 1.84 7.94 3.48 ;
        RECT  6.44 1.96 6.96 2.12 ;
        RECT  6.68 1.84 6.96 2.12 ;
        RECT  6.32 2.52 6.60 3.48 ;
        RECT  6.44 1.96 6.60 3.48 ;
        RECT  0.38 2.48 0.66 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 12.00 0.28 ;
        RECT  11.62 0.64 11.90 1.24 ;
        RECT  11.68 -0.28 11.84 1.24 ;
        RECT  11.54 -0.28 11.84 0.32 ;
        RECT  10.58 0.64 10.86 1.24 ;
        RECT  10.64 -0.28 10.80 1.24 ;
        RECT  8.75 0.88 9.10 1.16 ;
        RECT  8.75 -0.28 8.91 1.16 ;
        RECT  6.36 -0.28 6.64 0.68 ;
        RECT  0.38 -0.28 0.66 0.68 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  1.14 0.96 1.48 1.24 ;
        RECT  1.32 1.46 1.64 1.74 ;
        RECT  1.32 0.96 1.48 2.20 ;
        RECT  1.14 1.92 1.48 2.20 ;
        RECT  1.74 0.44 2.02 0.72 ;
        RECT  0.82 0.56 2.02 0.72 ;
        RECT  0.82 0.56 0.98 1.12 ;
        RECT  0.08 0.96 0.98 1.12 ;
        RECT  0.08 0.96 0.38 1.24 ;
        RECT  0.08 0.96 0.24 2.20 ;
        RECT  0.08 1.92 0.38 2.20 ;
        RECT  0.08 2.04 0.98 2.20 ;
        RECT  0.82 2.04 0.98 2.64 ;
        RECT  0.82 2.48 1.92 2.64 ;
        RECT  1.64 2.48 1.92 2.76 ;
        RECT  3.26 0.88 3.58 1.16 ;
        RECT  3.26 0.88 3.42 2.00 ;
        RECT  2.92 1.84 3.90 2.00 ;
        RECT  2.92 1.84 3.20 2.12 ;
        RECT  3.62 1.84 3.90 2.12 ;
        RECT  3.82 0.88 4.10 1.16 ;
        RECT  3.94 0.88 4.10 1.58 ;
        RECT  4.78 1.14 5.06 1.58 ;
        RECT  3.94 1.42 5.06 1.58 ;
        RECT  4.06 1.42 4.22 2.12 ;
        RECT  4.06 1.84 4.42 2.12 ;
        RECT  2.42 0.50 5.82 0.66 ;
        RECT  5.54 0.50 5.82 0.78 ;
        RECT  2.30 0.86 2.58 1.14 ;
        RECT  2.42 0.50 2.58 1.14 ;
        RECT  1.74 0.98 2.58 1.14 ;
        RECT  1.74 0.96 2.02 1.24 ;
        RECT  1.96 0.98 2.12 2.12 ;
        RECT  1.96 1.84 2.24 2.12 ;
        RECT  6.80 0.50 7.08 0.78 ;
        RECT  4.34 0.82 5.38 0.98 ;
        RECT  4.34 0.82 4.62 1.16 ;
        RECT  6.80 0.50 6.96 1.16 ;
        RECT  5.22 1.00 6.96 1.16 ;
        RECT  5.22 0.96 5.58 1.24 ;
        RECT  5.52 1.00 5.68 2.12 ;
        RECT  4.66 1.84 4.94 2.12 ;
        RECT  5.52 1.84 5.86 2.12 ;
        RECT  4.66 1.96 5.86 2.12 ;
        RECT  2.74 0.86 3.10 1.14 ;
        RECT  7.34 0.96 7.78 1.24 ;
        RECT  2.74 0.86 2.90 1.48 ;
        RECT  6.02 1.52 7.50 1.68 ;
        RECT  2.48 1.84 2.76 2.12 ;
        RECT  7.34 0.96 7.50 2.12 ;
        RECT  7.20 1.84 7.50 2.12 ;
        RECT  2.60 1.32 2.76 2.44 ;
        RECT  6.02 1.52 6.18 2.44 ;
        RECT  2.60 2.28 6.18 2.44 ;
        RECT  7.98 0.88 8.40 1.16 ;
        RECT  8.24 1.46 9.78 1.62 ;
        RECT  9.50 1.40 9.78 1.68 ;
        RECT  8.24 0.88 8.40 2.12 ;
        RECT  8.24 1.84 8.52 2.12 ;
        RECT  9.78 0.88 10.14 1.16 ;
        RECT  9.98 0.88 10.14 2.16 ;
        RECT  9.49 1.96 10.26 2.12 ;
        RECT  9.98 1.88 10.26 2.16 ;
        RECT  9.49 1.96 9.65 2.76 ;
        RECT  9.37 2.48 9.65 2.76 ;
    END
END DFFSRSSP4V1_0

MACRO DFFSRSSP2V1_0
    CLASS CORE ;
    FOREIGN DFFSRSSP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 22.23  LAYER ME1  ;
        ANTENNADIFFAREA 9.80  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.55  LAYER ME1  ;
        ANTENNAMAXAREACAR 40.62  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.22 1.46 11.52 1.74 ;
        RECT  11.10 1.84 11.38 2.44 ;
        RECT  11.22 0.64 11.38 2.44 ;
        RECT  11.10 0.64 11.38 1.24 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.40 0.70 1.76 ;
        END
    END D
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.66 1.40 8.08 1.68 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.40 1.16 1.76 ;
        END
    END CK
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.26 0.44 9.54 0.94 ;
        RECT  9.07 0.44 9.54 0.72 ;
        END
    END SB
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 11.60 0.28 ;
        RECT  11.14 -0.28 11.42 0.32 ;
        RECT  10.58 0.64 10.86 1.24 ;
        RECT  10.64 -0.28 10.80 1.24 ;
        RECT  8.75 0.88 9.10 1.16 ;
        RECT  8.75 -0.28 8.91 1.16 ;
        RECT  6.36 -0.28 6.64 0.68 ;
        RECT  0.38 -0.28 0.66 0.68 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 11.60 3.48 ;
        RECT  11.14 2.88 11.42 3.48 ;
        RECT  10.58 1.84 10.86 2.44 ;
        RECT  10.64 1.84 10.80 3.48 ;
        RECT  9.98 2.40 10.26 3.48 ;
        RECT  8.76 1.84 9.04 2.12 ;
        RECT  8.82 1.84 8.98 3.48 ;
        RECT  7.72 1.84 8.00 2.12 ;
        RECT  7.78 1.84 7.94 3.48 ;
        RECT  6.44 1.96 6.96 2.12 ;
        RECT  6.68 1.84 6.96 2.12 ;
        RECT  6.32 2.52 6.60 3.48 ;
        RECT  6.44 1.96 6.60 3.48 ;
        RECT  0.38 2.48 0.66 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  1.14 0.96 1.48 1.24 ;
        RECT  1.32 1.46 1.64 1.74 ;
        RECT  1.32 0.96 1.48 2.20 ;
        RECT  1.14 1.92 1.48 2.20 ;
        RECT  1.74 0.44 2.02 0.72 ;
        RECT  0.82 0.56 2.02 0.72 ;
        RECT  0.82 0.56 0.98 1.12 ;
        RECT  0.08 0.96 0.98 1.12 ;
        RECT  0.08 0.96 0.38 1.24 ;
        RECT  0.08 0.96 0.24 2.20 ;
        RECT  0.08 1.92 0.38 2.20 ;
        RECT  0.08 2.04 0.98 2.20 ;
        RECT  0.82 2.04 0.98 2.64 ;
        RECT  0.82 2.48 1.92 2.64 ;
        RECT  1.64 2.48 1.92 2.76 ;
        RECT  3.26 0.88 3.58 1.16 ;
        RECT  3.26 0.88 3.42 2.00 ;
        RECT  2.92 1.84 3.90 2.00 ;
        RECT  2.92 1.84 3.20 2.12 ;
        RECT  3.62 1.84 3.90 2.12 ;
        RECT  3.82 0.88 4.10 1.16 ;
        RECT  3.94 0.88 4.10 1.58 ;
        RECT  4.78 1.14 5.06 1.58 ;
        RECT  3.94 1.42 5.06 1.58 ;
        RECT  4.06 1.42 4.22 2.12 ;
        RECT  4.06 1.84 4.42 2.12 ;
        RECT  2.42 0.50 5.82 0.66 ;
        RECT  5.54 0.50 5.82 0.78 ;
        RECT  2.30 0.86 2.58 1.14 ;
        RECT  2.42 0.50 2.58 1.14 ;
        RECT  1.74 0.98 2.58 1.14 ;
        RECT  1.74 0.96 2.02 1.24 ;
        RECT  1.96 0.98 2.12 2.12 ;
        RECT  1.96 1.84 2.24 2.12 ;
        RECT  6.80 0.50 7.08 0.78 ;
        RECT  4.34 0.82 5.38 0.98 ;
        RECT  4.34 0.82 4.62 1.16 ;
        RECT  6.80 0.50 6.96 1.16 ;
        RECT  5.22 1.00 6.96 1.16 ;
        RECT  5.22 0.96 5.58 1.24 ;
        RECT  5.52 1.00 5.68 2.12 ;
        RECT  4.66 1.84 4.94 2.12 ;
        RECT  5.52 1.84 5.86 2.12 ;
        RECT  4.66 1.96 5.86 2.12 ;
        RECT  2.74 0.86 3.10 1.14 ;
        RECT  7.34 0.96 7.78 1.24 ;
        RECT  2.74 0.86 2.90 1.48 ;
        RECT  6.02 1.52 7.50 1.68 ;
        RECT  2.48 1.84 2.76 2.12 ;
        RECT  7.34 0.96 7.50 2.12 ;
        RECT  7.20 1.84 7.50 2.12 ;
        RECT  2.60 1.32 2.76 2.44 ;
        RECT  6.02 1.52 6.18 2.44 ;
        RECT  2.60 2.28 6.18 2.44 ;
        RECT  7.98 0.88 8.40 1.16 ;
        RECT  8.24 1.46 9.78 1.62 ;
        RECT  9.50 1.40 9.78 1.68 ;
        RECT  8.24 0.88 8.40 2.12 ;
        RECT  8.24 1.84 8.52 2.12 ;
        RECT  9.78 0.88 10.14 1.16 ;
        RECT  9.98 0.88 10.14 2.16 ;
        RECT  9.49 1.96 10.26 2.12 ;
        RECT  9.98 1.88 10.26 2.16 ;
        RECT  9.49 1.96 9.65 2.76 ;
        RECT  9.37 2.48 9.65 2.76 ;
    END
END DFFSRSSP2V1_0

MACRO DFFSRSSP1V1_0
    CLASS CORE ;
    FOREIGN DFFSRSSP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 21.68  LAYER ME1  ;
        ANTENNADIFFAREA 9.36  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.47  LAYER ME1  ;
        ANTENNAMAXAREACAR 46.09  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.22 1.46 11.52 1.74 ;
        RECT  11.10 1.84 11.38 2.12 ;
        RECT  11.22 0.96 11.38 2.12 ;
        RECT  11.10 0.96 11.38 1.24 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.40 0.70 1.76 ;
        END
    END D
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.66 1.40 8.08 1.68 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.40 1.16 1.76 ;
        END
    END CK
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.26 0.44 9.54 0.94 ;
        RECT  9.07 0.44 9.54 0.72 ;
        END
    END SB
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 11.60 3.48 ;
        RECT  11.14 2.88 11.42 3.48 ;
        RECT  10.58 1.84 10.86 2.12 ;
        RECT  10.64 1.84 10.80 3.48 ;
        RECT  9.98 2.40 10.26 3.48 ;
        RECT  8.76 1.84 9.04 2.12 ;
        RECT  8.82 1.84 8.98 3.48 ;
        RECT  7.72 1.84 8.00 2.12 ;
        RECT  7.78 1.84 7.94 3.48 ;
        RECT  6.44 1.96 6.96 2.12 ;
        RECT  6.68 1.84 6.96 2.12 ;
        RECT  6.32 2.52 6.60 3.48 ;
        RECT  6.44 1.96 6.60 3.48 ;
        RECT  0.38 2.48 0.66 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 11.60 0.28 ;
        RECT  11.14 -0.28 11.42 0.32 ;
        RECT  10.58 0.96 10.86 1.24 ;
        RECT  10.64 -0.28 10.80 1.24 ;
        RECT  8.75 0.88 9.10 1.16 ;
        RECT  8.75 -0.28 8.91 1.16 ;
        RECT  6.36 -0.28 6.64 0.68 ;
        RECT  0.38 -0.28 0.66 0.68 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  1.14 0.96 1.48 1.24 ;
        RECT  1.32 1.46 1.64 1.74 ;
        RECT  1.32 0.96 1.48 2.20 ;
        RECT  1.14 1.92 1.48 2.20 ;
        RECT  1.74 0.44 2.02 0.72 ;
        RECT  0.82 0.56 2.02 0.72 ;
        RECT  0.82 0.56 0.98 1.12 ;
        RECT  0.08 0.96 0.98 1.12 ;
        RECT  0.08 0.96 0.38 1.24 ;
        RECT  0.08 0.96 0.24 2.20 ;
        RECT  0.08 1.92 0.38 2.20 ;
        RECT  0.08 2.04 0.98 2.20 ;
        RECT  0.82 2.04 0.98 2.64 ;
        RECT  0.82 2.48 1.92 2.64 ;
        RECT  1.64 2.48 1.92 2.76 ;
        RECT  3.26 0.88 3.58 1.16 ;
        RECT  3.26 0.88 3.42 2.00 ;
        RECT  2.92 1.84 3.90 2.00 ;
        RECT  2.92 1.84 3.20 2.12 ;
        RECT  3.62 1.84 3.90 2.12 ;
        RECT  3.82 0.88 4.10 1.16 ;
        RECT  3.94 0.88 4.10 1.58 ;
        RECT  4.78 1.14 5.06 1.58 ;
        RECT  3.94 1.42 5.06 1.58 ;
        RECT  4.06 1.42 4.22 2.12 ;
        RECT  4.06 1.84 4.42 2.12 ;
        RECT  2.42 0.50 5.82 0.66 ;
        RECT  5.54 0.50 5.82 0.78 ;
        RECT  2.30 0.86 2.58 1.14 ;
        RECT  2.42 0.50 2.58 1.14 ;
        RECT  1.74 0.98 2.58 1.14 ;
        RECT  1.74 0.96 2.02 1.24 ;
        RECT  1.96 0.98 2.12 2.12 ;
        RECT  1.96 1.84 2.24 2.12 ;
        RECT  6.80 0.50 7.08 0.78 ;
        RECT  4.34 0.82 5.38 0.98 ;
        RECT  4.34 0.82 4.62 1.16 ;
        RECT  6.80 0.50 6.96 1.16 ;
        RECT  5.22 1.00 6.96 1.16 ;
        RECT  5.22 0.96 5.58 1.24 ;
        RECT  5.52 1.00 5.68 2.12 ;
        RECT  4.66 1.84 4.94 2.12 ;
        RECT  5.52 1.84 5.86 2.12 ;
        RECT  4.66 1.96 5.86 2.12 ;
        RECT  2.74 0.86 3.10 1.14 ;
        RECT  7.34 0.96 7.78 1.24 ;
        RECT  2.74 0.86 2.90 1.48 ;
        RECT  6.02 1.52 7.50 1.68 ;
        RECT  2.48 1.84 2.76 2.12 ;
        RECT  7.34 0.96 7.50 2.12 ;
        RECT  7.20 1.84 7.50 2.12 ;
        RECT  2.60 1.32 2.76 2.44 ;
        RECT  6.02 1.52 6.18 2.44 ;
        RECT  2.60 2.28 6.18 2.44 ;
        RECT  7.98 0.88 8.40 1.16 ;
        RECT  8.24 1.46 9.78 1.62 ;
        RECT  9.50 1.40 9.78 1.68 ;
        RECT  8.24 0.88 8.40 2.12 ;
        RECT  8.24 1.84 8.52 2.12 ;
        RECT  9.78 0.88 10.14 1.16 ;
        RECT  9.98 0.88 10.14 2.16 ;
        RECT  9.49 1.96 10.26 2.12 ;
        RECT  9.98 1.88 10.26 2.16 ;
        RECT  9.49 1.96 9.65 2.76 ;
        RECT  9.37 2.48 9.65 2.76 ;
    END
END DFFSRSSP1V1_0

MACRO DFFSRSP8V1_0
    CLASS CORE ;
    FOREIGN DFFSRSP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.42 2.28 6.80 2.56 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.88 1.40 1.20 1.76 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.40 0.72 1.76 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 22.90  LAYER ME1  ;
        ANTENNADIFFAREA 10.84  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.98  LAYER ME1  ;
        ANTENNAMAXAREACAR 23.39  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.50 1.90 10.78 2.50 ;
        RECT  10.50 0.64 10.78 1.24 ;
        RECT  10.50 0.64 10.66 2.50 ;
        RECT  9.26 1.52 10.66 1.68 ;
        RECT  9.46 1.90 9.74 2.50 ;
        RECT  9.46 0.64 9.74 1.24 ;
        RECT  9.46 0.64 9.62 2.50 ;
        RECT  9.26 1.46 9.62 1.74 ;
        END
    END Q
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 11.60 0.28 ;
        RECT  11.08 -0.28 11.42 0.32 ;
        RECT  11.02 0.64 11.30 1.24 ;
        RECT  11.08 -0.28 11.24 1.24 ;
        RECT  9.98 0.64 10.26 1.24 ;
        RECT  10.04 -0.28 10.20 1.24 ;
        RECT  8.94 0.64 9.22 1.24 ;
        RECT  9.00 -0.28 9.16 1.24 ;
        RECT  7.94 0.88 8.22 1.16 ;
        RECT  8.00 -0.28 8.16 1.16 ;
        RECT  4.96 -0.28 5.24 0.72 ;
        RECT  0.38 -0.28 0.66 0.68 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 11.60 3.48 ;
        RECT  11.08 2.88 11.42 3.48 ;
        RECT  11.02 1.90 11.30 2.50 ;
        RECT  11.08 1.90 11.24 3.48 ;
        RECT  9.98 1.90 10.26 2.50 ;
        RECT  10.04 1.90 10.20 3.48 ;
        RECT  8.94 1.90 9.22 2.50 ;
        RECT  9.00 1.90 9.16 3.48 ;
        RECT  7.94 1.84 8.22 2.12 ;
        RECT  8.00 1.84 8.16 3.48 ;
        RECT  7.10 1.84 7.26 3.48 ;
        RECT  6.90 1.84 7.26 2.12 ;
        RECT  6.06 1.84 6.22 3.48 ;
        RECT  5.86 1.84 6.22 2.12 ;
        RECT  0.38 2.48 0.66 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  1.14 0.96 1.52 1.24 ;
        RECT  1.36 1.46 1.64 1.74 ;
        RECT  1.36 0.96 1.52 2.20 ;
        RECT  1.14 1.92 1.52 2.20 ;
        RECT  1.74 0.44 2.02 0.72 ;
        RECT  0.82 0.56 2.02 0.72 ;
        RECT  0.82 0.56 0.98 1.12 ;
        RECT  0.08 0.96 0.98 1.12 ;
        RECT  0.08 0.96 0.38 1.24 ;
        RECT  0.08 0.96 0.24 2.20 ;
        RECT  0.08 1.92 0.38 2.20 ;
        RECT  0.08 2.04 0.98 2.20 ;
        RECT  0.82 2.04 0.98 2.64 ;
        RECT  0.82 2.48 2.02 2.64 ;
        RECT  1.74 2.48 2.02 2.76 ;
        RECT  3.34 0.88 3.62 1.16 ;
        RECT  3.34 0.88 3.50 2.12 ;
        RECT  3.12 1.84 3.50 2.12 ;
        RECT  3.82 1.84 4.10 2.12 ;
        RECT  3.12 1.96 4.10 2.12 ;
        RECT  4.52 0.44 4.80 0.72 ;
        RECT  3.98 0.56 4.80 0.72 ;
        RECT  3.86 0.88 4.14 1.16 ;
        RECT  3.98 0.56 4.14 1.68 ;
        RECT  3.98 1.52 4.42 1.68 ;
        RECT  4.26 1.52 4.42 2.12 ;
        RECT  4.26 1.84 4.62 2.12 ;
        RECT  2.30 0.87 2.58 1.15 ;
        RECT  1.74 0.99 2.58 1.15 ;
        RECT  1.74 0.96 2.02 1.24 ;
        RECT  1.86 0.96 2.02 2.12 ;
        RECT  1.86 1.84 2.14 2.12 ;
        RECT  1.86 1.96 2.44 2.12 ;
        RECT  2.28 1.96 2.44 2.76 ;
        RECT  5.62 2.42 5.90 2.76 ;
        RECT  2.28 2.60 5.90 2.76 ;
        RECT  5.82 0.50 6.10 0.78 ;
        RECT  4.38 0.88 4.66 1.20 ;
        RECT  5.00 0.92 5.28 1.20 ;
        RECT  5.82 0.50 5.98 1.20 ;
        RECT  4.38 1.04 5.98 1.20 ;
        RECT  4.78 1.04 4.94 2.12 ;
        RECT  4.78 1.84 5.14 2.12 ;
        RECT  2.80 0.87 3.10 1.15 ;
        RECT  6.48 0.92 6.76 1.20 ;
        RECT  5.30 1.52 6.64 1.68 ;
        RECT  6.48 0.92 6.64 2.12 ;
        RECT  2.68 1.84 2.96 2.12 ;
        RECT  6.38 1.84 6.66 2.12 ;
        RECT  2.80 0.87 2.96 2.44 ;
        RECT  5.30 1.52 5.46 2.44 ;
        RECT  2.80 2.28 5.46 2.44 ;
        RECT  7.04 0.88 7.32 1.16 ;
        RECT  7.04 1.00 7.58 1.16 ;
        RECT  7.42 1.46 8.42 1.62 ;
        RECT  8.14 1.40 8.42 1.68 ;
        RECT  7.42 1.00 7.58 2.12 ;
        RECT  7.42 1.84 7.70 2.12 ;
        RECT  8.46 0.88 8.74 1.16 ;
        RECT  8.46 1.84 8.74 2.12 ;
        RECT  8.58 0.88 8.74 2.76 ;
        RECT  8.49 2.48 8.77 2.76 ;
    END
END DFFSRSP8V1_0

MACRO DFFSRSP4V1_0
    CLASS CORE ;
    FOREIGN DFFSRSP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 20.51  LAYER ME1  ;
        ANTENNADIFFAREA 9.02  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.69  LAYER ME1  ;
        ANTENNAMAXAREACAR 29.67  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.46 1.90 9.74 2.50 ;
        RECT  9.46 0.64 9.74 1.24 ;
        RECT  9.46 0.64 9.62 2.50 ;
        RECT  9.26 1.46 9.62 1.74 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.40 0.72 1.76 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.88 1.40 1.20 1.76 ;
        END
    END CK
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.42 2.28 6.80 2.56 ;
        END
    END RB
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 10.40 3.48 ;
        RECT  9.98 1.90 10.26 2.50 ;
        RECT  9.94 2.88 10.22 3.48 ;
        RECT  10.04 1.90 10.20 3.48 ;
        RECT  8.94 1.90 9.22 2.50 ;
        RECT  9.00 1.90 9.16 3.48 ;
        RECT  7.94 1.84 8.22 2.12 ;
        RECT  8.00 1.84 8.16 3.48 ;
        RECT  7.10 1.84 7.26 3.48 ;
        RECT  6.90 1.84 7.26 2.12 ;
        RECT  6.06 1.84 6.22 3.48 ;
        RECT  5.86 1.84 6.22 2.12 ;
        RECT  0.38 2.48 0.66 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 10.40 0.28 ;
        RECT  9.98 0.64 10.26 1.24 ;
        RECT  9.94 -0.28 10.22 0.32 ;
        RECT  10.04 -0.28 10.20 1.24 ;
        RECT  8.94 0.64 9.22 1.24 ;
        RECT  9.00 -0.28 9.16 1.24 ;
        RECT  7.94 0.88 8.22 1.16 ;
        RECT  8.00 -0.28 8.16 1.16 ;
        RECT  4.96 -0.28 5.24 0.72 ;
        RECT  0.38 -0.28 0.66 0.68 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  1.14 0.96 1.52 1.24 ;
        RECT  1.36 1.46 1.64 1.74 ;
        RECT  1.36 0.96 1.52 2.20 ;
        RECT  1.14 1.92 1.52 2.20 ;
        RECT  1.74 0.44 2.02 0.72 ;
        RECT  0.82 0.56 2.02 0.72 ;
        RECT  0.82 0.56 0.98 1.12 ;
        RECT  0.08 0.96 0.98 1.12 ;
        RECT  0.08 0.96 0.38 1.24 ;
        RECT  0.08 0.96 0.24 2.20 ;
        RECT  0.08 1.92 0.38 2.20 ;
        RECT  0.08 2.04 0.98 2.20 ;
        RECT  0.82 2.04 0.98 2.64 ;
        RECT  0.82 2.48 2.02 2.64 ;
        RECT  1.74 2.48 2.02 2.76 ;
        RECT  3.34 0.88 3.62 1.16 ;
        RECT  3.34 0.88 3.50 2.12 ;
        RECT  3.12 1.84 3.50 2.12 ;
        RECT  3.82 1.84 4.10 2.12 ;
        RECT  3.12 1.96 4.10 2.12 ;
        RECT  4.52 0.44 4.80 0.72 ;
        RECT  3.98 0.56 4.80 0.72 ;
        RECT  3.86 0.88 4.14 1.16 ;
        RECT  3.98 0.56 4.14 1.68 ;
        RECT  3.98 1.52 4.42 1.68 ;
        RECT  4.26 1.52 4.42 2.12 ;
        RECT  4.26 1.84 4.62 2.12 ;
        RECT  2.30 0.87 2.58 1.15 ;
        RECT  1.74 0.99 2.58 1.15 ;
        RECT  1.74 0.96 2.02 1.24 ;
        RECT  1.86 0.96 2.02 2.12 ;
        RECT  1.86 1.84 2.14 2.12 ;
        RECT  1.86 1.96 2.44 2.12 ;
        RECT  2.28 1.96 2.44 2.76 ;
        RECT  5.62 2.42 5.90 2.76 ;
        RECT  2.28 2.60 5.90 2.76 ;
        RECT  5.82 0.50 6.10 0.78 ;
        RECT  4.38 0.88 4.66 1.20 ;
        RECT  5.00 0.92 5.28 1.20 ;
        RECT  5.82 0.50 5.98 1.20 ;
        RECT  4.38 1.04 5.98 1.20 ;
        RECT  4.78 1.04 4.94 2.12 ;
        RECT  4.78 1.84 5.14 2.12 ;
        RECT  2.80 0.87 3.10 1.15 ;
        RECT  6.48 0.92 6.76 1.20 ;
        RECT  5.30 1.52 6.64 1.68 ;
        RECT  6.48 0.92 6.64 2.12 ;
        RECT  2.68 1.84 2.96 2.12 ;
        RECT  6.38 1.84 6.66 2.12 ;
        RECT  2.80 0.87 2.96 2.44 ;
        RECT  5.30 1.52 5.46 2.44 ;
        RECT  2.80 2.28 5.46 2.44 ;
        RECT  7.04 0.88 7.32 1.16 ;
        RECT  7.04 1.00 7.58 1.16 ;
        RECT  7.42 1.46 8.42 1.62 ;
        RECT  8.14 1.40 8.42 1.68 ;
        RECT  7.42 1.00 7.58 2.12 ;
        RECT  7.42 1.84 7.70 2.12 ;
        RECT  8.46 0.88 8.74 1.16 ;
        RECT  8.46 1.84 8.74 2.12 ;
        RECT  8.58 0.88 8.74 2.76 ;
        RECT  8.49 2.48 8.77 2.76 ;
    END
END DFFSRSP4V1_0

MACRO DFFSRSP2V1_0
    CLASS CORE ;
    FOREIGN DFFSRSP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.42 2.28 6.80 2.56 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.88 1.40 1.20 1.76 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.40 0.72 1.76 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 19.62  LAYER ME1  ;
        ANTENNADIFFAREA 8.41  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.55  LAYER ME1  ;
        ANTENNAMAXAREACAR 35.85  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.46 1.90 9.74 2.50 ;
        RECT  9.46 0.64 9.74 1.24 ;
        RECT  9.46 0.64 9.62 2.50 ;
        RECT  9.26 1.46 9.62 1.74 ;
        END
    END Q
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 10.00 0.28 ;
        RECT  9.54 -0.28 9.82 0.32 ;
        RECT  8.94 0.64 9.22 1.24 ;
        RECT  9.00 -0.28 9.16 1.24 ;
        RECT  7.94 0.88 8.22 1.16 ;
        RECT  8.00 -0.28 8.16 1.16 ;
        RECT  4.96 -0.28 5.24 0.72 ;
        RECT  0.38 -0.28 0.66 0.68 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 10.00 3.48 ;
        RECT  9.54 2.88 9.82 3.48 ;
        RECT  8.94 1.90 9.22 2.50 ;
        RECT  9.00 1.90 9.16 3.48 ;
        RECT  7.94 1.84 8.22 2.12 ;
        RECT  8.00 1.84 8.16 3.48 ;
        RECT  7.10 1.84 7.26 3.48 ;
        RECT  6.90 1.84 7.26 2.12 ;
        RECT  6.06 1.84 6.22 3.48 ;
        RECT  5.86 1.84 6.22 2.12 ;
        RECT  0.38 2.48 0.66 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  1.14 0.96 1.52 1.24 ;
        RECT  1.36 1.46 1.64 1.74 ;
        RECT  1.36 0.96 1.52 2.20 ;
        RECT  1.14 1.92 1.52 2.20 ;
        RECT  1.74 0.44 2.02 0.72 ;
        RECT  0.82 0.56 2.02 0.72 ;
        RECT  0.82 0.56 0.98 1.12 ;
        RECT  0.08 0.96 0.98 1.12 ;
        RECT  0.08 0.96 0.38 1.24 ;
        RECT  0.08 0.96 0.24 2.20 ;
        RECT  0.08 1.92 0.38 2.20 ;
        RECT  0.08 2.04 0.98 2.20 ;
        RECT  0.82 2.04 0.98 2.64 ;
        RECT  0.82 2.48 2.02 2.64 ;
        RECT  1.74 2.48 2.02 2.76 ;
        RECT  3.34 0.88 3.62 1.16 ;
        RECT  3.34 0.88 3.50 2.12 ;
        RECT  3.12 1.84 3.50 2.12 ;
        RECT  3.82 1.84 4.10 2.12 ;
        RECT  3.12 1.96 4.10 2.12 ;
        RECT  4.52 0.44 4.80 0.72 ;
        RECT  3.98 0.56 4.80 0.72 ;
        RECT  3.86 0.88 4.14 1.16 ;
        RECT  3.98 0.56 4.14 1.68 ;
        RECT  3.98 1.52 4.42 1.68 ;
        RECT  4.26 1.52 4.42 2.12 ;
        RECT  4.26 1.84 4.62 2.12 ;
        RECT  2.30 0.87 2.58 1.15 ;
        RECT  1.74 0.99 2.58 1.15 ;
        RECT  1.74 0.96 2.02 1.24 ;
        RECT  1.86 0.96 2.02 2.12 ;
        RECT  1.86 1.84 2.14 2.12 ;
        RECT  1.86 1.96 2.44 2.12 ;
        RECT  2.28 1.96 2.44 2.76 ;
        RECT  5.62 2.42 5.90 2.76 ;
        RECT  2.28 2.60 5.90 2.76 ;
        RECT  5.82 0.50 6.10 0.78 ;
        RECT  4.38 0.88 4.66 1.20 ;
        RECT  5.00 0.92 5.28 1.20 ;
        RECT  5.82 0.50 5.98 1.20 ;
        RECT  4.38 1.04 5.98 1.20 ;
        RECT  4.78 1.04 4.94 2.12 ;
        RECT  4.78 1.84 5.14 2.12 ;
        RECT  2.80 0.87 3.10 1.15 ;
        RECT  6.48 0.92 6.76 1.20 ;
        RECT  5.30 1.52 6.64 1.68 ;
        RECT  6.48 0.92 6.64 2.12 ;
        RECT  2.68 1.84 2.96 2.12 ;
        RECT  6.38 1.84 6.66 2.12 ;
        RECT  2.80 0.87 2.96 2.44 ;
        RECT  5.30 1.52 5.46 2.44 ;
        RECT  2.80 2.28 5.46 2.44 ;
        RECT  7.04 0.88 7.32 1.16 ;
        RECT  7.04 1.00 7.58 1.16 ;
        RECT  7.42 1.46 8.42 1.62 ;
        RECT  8.14 1.40 8.42 1.68 ;
        RECT  7.42 1.00 7.58 2.12 ;
        RECT  7.42 1.84 7.70 2.12 ;
        RECT  8.46 0.88 8.74 1.16 ;
        RECT  8.46 1.84 8.74 2.12 ;
        RECT  8.58 0.88 8.74 2.76 ;
        RECT  8.49 2.48 8.77 2.76 ;
    END
END DFFSRSP2V1_0

MACRO DFFSRSP1V1_0
    CLASS CORE ;
    FOREIGN DFFSRSP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 19.03  LAYER ME1  ;
        ANTENNADIFFAREA 7.98  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.47  LAYER ME1  ;
        ANTENNAMAXAREACAR 40.45  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.46 1.90 9.74 2.18 ;
        RECT  9.46 0.88 9.74 1.16 ;
        RECT  9.46 0.88 9.62 2.18 ;
        RECT  9.26 1.46 9.62 1.74 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.40 0.72 1.76 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.88 1.40 1.20 1.76 ;
        END
    END CK
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.42 2.28 6.80 2.56 ;
        END
    END RB
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 10.00 0.28 ;
        RECT  9.54 -0.28 9.82 0.32 ;
        RECT  8.94 0.88 9.22 1.16 ;
        RECT  9.00 -0.28 9.16 1.16 ;
        RECT  7.94 0.88 8.22 1.16 ;
        RECT  8.00 -0.28 8.16 1.16 ;
        RECT  4.96 -0.28 5.24 0.72 ;
        RECT  0.38 -0.28 0.66 0.68 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 10.00 3.48 ;
        RECT  9.54 2.88 9.82 3.48 ;
        RECT  8.94 1.90 9.22 2.18 ;
        RECT  9.00 1.90 9.16 3.48 ;
        RECT  7.94 1.84 8.22 2.12 ;
        RECT  8.00 1.84 8.16 3.48 ;
        RECT  7.10 1.84 7.26 3.48 ;
        RECT  6.90 1.84 7.26 2.12 ;
        RECT  6.06 1.84 6.22 3.48 ;
        RECT  5.86 1.84 6.22 2.12 ;
        RECT  0.38 2.48 0.66 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  1.14 0.96 1.52 1.24 ;
        RECT  1.36 1.46 1.64 1.74 ;
        RECT  1.36 0.96 1.52 2.20 ;
        RECT  1.14 1.92 1.52 2.20 ;
        RECT  1.74 0.44 2.02 0.72 ;
        RECT  0.82 0.56 2.02 0.72 ;
        RECT  0.82 0.56 0.98 1.12 ;
        RECT  0.08 0.96 0.98 1.12 ;
        RECT  0.08 0.96 0.38 1.24 ;
        RECT  0.08 0.96 0.24 2.20 ;
        RECT  0.08 1.92 0.38 2.20 ;
        RECT  0.08 2.04 0.98 2.20 ;
        RECT  0.82 2.04 0.98 2.64 ;
        RECT  0.82 2.48 2.02 2.64 ;
        RECT  1.74 2.48 2.02 2.76 ;
        RECT  3.34 0.88 3.62 1.16 ;
        RECT  3.34 0.88 3.50 2.12 ;
        RECT  3.12 1.84 3.50 2.12 ;
        RECT  3.82 1.84 4.10 2.12 ;
        RECT  3.12 1.96 4.10 2.12 ;
        RECT  4.52 0.44 4.80 0.72 ;
        RECT  3.98 0.56 4.80 0.72 ;
        RECT  3.86 0.88 4.14 1.16 ;
        RECT  3.98 0.56 4.14 1.68 ;
        RECT  3.98 1.52 4.42 1.68 ;
        RECT  4.26 1.52 4.42 2.12 ;
        RECT  4.26 1.84 4.62 2.12 ;
        RECT  2.30 0.87 2.58 1.15 ;
        RECT  1.74 0.99 2.58 1.15 ;
        RECT  1.74 0.96 2.02 1.24 ;
        RECT  1.86 0.96 2.02 2.12 ;
        RECT  1.86 1.84 2.14 2.12 ;
        RECT  1.86 1.96 2.44 2.12 ;
        RECT  2.28 1.96 2.44 2.76 ;
        RECT  5.62 2.42 5.90 2.76 ;
        RECT  2.28 2.60 5.90 2.76 ;
        RECT  5.82 0.50 6.10 0.78 ;
        RECT  4.38 0.88 4.66 1.20 ;
        RECT  5.00 0.92 5.28 1.20 ;
        RECT  5.82 0.50 5.98 1.20 ;
        RECT  4.38 1.04 5.98 1.20 ;
        RECT  4.78 1.04 4.94 2.12 ;
        RECT  4.78 1.84 5.14 2.12 ;
        RECT  2.80 0.87 3.10 1.15 ;
        RECT  6.48 0.92 6.76 1.20 ;
        RECT  5.30 1.52 6.64 1.68 ;
        RECT  6.48 0.92 6.64 2.12 ;
        RECT  2.68 1.84 2.96 2.12 ;
        RECT  6.38 1.84 6.66 2.12 ;
        RECT  2.80 0.87 2.96 2.44 ;
        RECT  5.30 1.52 5.46 2.44 ;
        RECT  2.80 2.28 5.46 2.44 ;
        RECT  7.04 0.88 7.32 1.16 ;
        RECT  7.04 1.00 7.58 1.16 ;
        RECT  7.42 1.46 8.42 1.62 ;
        RECT  8.14 1.40 8.42 1.68 ;
        RECT  7.42 1.00 7.58 2.12 ;
        RECT  7.42 1.84 7.70 2.12 ;
        RECT  8.46 0.88 8.74 1.16 ;
        RECT  8.46 1.84 8.74 2.12 ;
        RECT  8.58 0.88 8.74 2.76 ;
        RECT  8.49 2.48 8.77 2.76 ;
    END
END DFFSRSP1V1_0

MACRO DFFDZSP8V1_1
    CLASS CORE ;
    FOREIGN DFFDZSP8V1_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 24.64  LAYER ME1  ;
        ANTENNADIFFAREA 12.66  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.62  LAYER ME1  ;
        ANTENNAMAXAREACAR 15.19  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.97 1.84 13.25 2.12 ;
        RECT  12.97 0.96 13.25 1.24 ;
        RECT  12.97 0.96 13.13 2.12 ;
        RECT  12.05 1.52 13.13 1.68 ;
        RECT  12.05 1.46 12.34 1.74 ;
        RECT  11.93 1.84 12.21 2.12 ;
        RECT  12.05 0.96 12.21 2.12 ;
        RECT  11.93 0.96 12.21 1.24 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 24.64  LAYER ME1  ;
        ANTENNADIFFAREA 12.66  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.62  LAYER ME1  ;
        ANTENNAMAXAREACAR 15.19  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.89 1.84 11.17 2.12 ;
        RECT  10.89 0.96 11.17 1.24 ;
        RECT  10.89 0.96 11.05 2.12 ;
        RECT  9.97 1.52 11.05 1.68 ;
        RECT  9.97 1.46 10.34 1.74 ;
        RECT  9.85 1.84 10.13 2.12 ;
        RECT  9.97 0.96 10.13 2.12 ;
        RECT  9.85 0.96 10.13 1.24 ;
        END
    END QB
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.92  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 13.64  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.07 1.46 2.32 1.74 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.81 2.23 2.25 ;
        RECT  1.95 0.81 2.23 1.09 ;
        END
    END TD
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END SEL
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.86 1.46 3.37 1.74 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.24  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 18.44  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.81 1.19 2.25 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  0.91 0.81 1.19 1.09 ;
        END
    END D
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 14.00 3.48 ;
        RECT  13.54 2.88 13.82 3.48 ;
        RECT  13.49 2.16 13.77 2.44 ;
        RECT  13.55 2.16 13.71 3.48 ;
        RECT  12.45 2.16 12.73 2.44 ;
        RECT  12.51 2.16 12.67 3.48 ;
        RECT  11.41 2.16 11.69 2.44 ;
        RECT  11.47 2.16 11.63 3.48 ;
        RECT  10.37 2.16 10.65 2.44 ;
        RECT  10.43 2.16 10.59 3.48 ;
        RECT  9.33 1.84 9.61 2.12 ;
        RECT  9.39 1.84 9.55 3.48 ;
        RECT  8.33 2.62 8.61 3.48 ;
        RECT  5.77 1.92 6.05 2.20 ;
        RECT  5.83 1.92 5.99 3.48 ;
        RECT  2.95 2.62 3.23 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 14.00 0.28 ;
        RECT  13.54 -0.28 13.82 0.32 ;
        RECT  13.49 0.64 13.77 0.92 ;
        RECT  13.55 -0.28 13.71 0.92 ;
        RECT  12.45 0.64 12.73 0.92 ;
        RECT  12.51 -0.28 12.67 0.92 ;
        RECT  11.41 0.64 11.69 0.92 ;
        RECT  11.47 -0.28 11.63 0.92 ;
        RECT  10.37 0.64 10.65 0.92 ;
        RECT  10.43 -0.28 10.59 0.92 ;
        RECT  9.33 0.64 9.61 0.92 ;
        RECT  9.39 -0.28 9.55 0.92 ;
        RECT  8.33 0.96 8.61 1.24 ;
        RECT  8.43 -0.28 8.59 1.24 ;
        RECT  5.59 0.72 5.87 1.00 ;
        RECT  5.65 -0.28 5.81 1.00 ;
        RECT  2.95 0.87 3.23 1.15 ;
        RECT  3.01 -0.28 3.17 1.15 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  1.55 1.97 1.71 2.58 ;
        RECT  2.39 2.30 2.67 2.58 ;
        RECT  1.55 2.42 2.67 2.58 ;
        RECT  3.47 0.87 3.77 1.15 ;
        RECT  3.61 1.25 3.89 1.53 ;
        RECT  3.61 0.87 3.77 2.14 ;
        RECT  3.49 1.86 3.77 2.14 ;
        RECT  3.97 0.72 4.25 1.00 ;
        RECT  2.43 0.87 2.71 1.15 ;
        RECT  2.54 0.87 2.70 2.14 ;
        RECT  4.05 0.72 4.21 2.20 ;
        RECT  2.43 1.86 2.71 2.14 ;
        RECT  2.43 1.98 3.07 2.14 ;
        RECT  3.97 1.92 4.25 2.20 ;
        RECT  2.91 1.98 3.07 2.46 ;
        RECT  3.97 1.92 4.13 2.46 ;
        RECT  2.91 2.30 4.13 2.46 ;
        RECT  5.05 0.72 5.35 1.00 ;
        RECT  5.05 0.72 5.21 2.20 ;
        RECT  5.01 1.92 5.29 2.20 ;
        RECT  4.49 0.72 4.77 1.00 ;
        RECT  5.85 1.48 6.13 1.76 ;
        RECT  5.45 1.60 6.13 1.76 ;
        RECT  4.55 0.72 4.71 2.20 ;
        RECT  4.49 1.92 4.77 2.20 ;
        RECT  4.61 1.92 4.77 2.52 ;
        RECT  5.45 1.60 5.61 2.52 ;
        RECT  4.61 2.36 5.61 2.52 ;
        RECT  6.11 0.72 6.45 1.00 ;
        RECT  5.37 1.16 6.45 1.32 ;
        RECT  5.37 1.16 5.65 1.44 ;
        RECT  6.29 0.72 6.45 2.20 ;
        RECT  6.29 1.92 6.57 2.20 ;
        RECT  6.79 0.44 8.27 0.60 ;
        RECT  7.99 0.44 8.27 0.80 ;
        RECT  6.67 0.76 6.95 1.04 ;
        RECT  6.79 0.44 6.95 2.20 ;
        RECT  6.79 1.92 7.09 2.20 ;
        RECT  7.81 0.96 8.09 1.24 ;
        RECT  7.81 1.46 8.78 1.62 ;
        RECT  8.50 1.40 8.78 1.68 ;
        RECT  7.81 0.96 7.97 2.12 ;
        RECT  7.81 1.84 8.09 2.12 ;
        RECT  7.19 0.76 7.49 1.04 ;
        RECT  8.85 0.96 9.13 1.24 ;
        RECT  8.85 1.84 9.13 2.12 ;
        RECT  7.33 0.76 7.49 2.20 ;
        RECT  7.45 1.92 7.61 2.44 ;
        RECT  8.94 0.96 9.10 2.70 ;
        RECT  7.45 2.28 9.10 2.44 ;
        RECT  8.94 2.42 9.23 2.70 ;
    END
END DFFDZSP8V1_1

MACRO DFFDZSP8V1_0
    CLASS CORE ;
    FOREIGN DFFDZSP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 27.59  LAYER ME1  ;
        ANTENNADIFFAREA 13.79  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.92  LAYER ME1  ;
        ANTENNAMAXAREACAR 14.33  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.12 1.84 14.42 2.12 ;
        RECT  14.12 0.96 14.42 1.24 ;
        RECT  14.12 0.96 14.28 2.12 ;
        RECT  13.22 1.52 14.28 1.68 ;
        RECT  13.10 1.84 13.38 2.12 ;
        RECT  13.22 0.96 13.38 2.12 ;
        RECT  13.10 0.96 13.38 1.24 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 27.59  LAYER ME1  ;
        ANTENNADIFFAREA 13.99  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.92  LAYER ME1  ;
        ANTENNAMAXAREACAR 14.33  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.06 1.84 12.34 2.12 ;
        RECT  12.06 0.96 12.34 1.24 ;
        RECT  12.06 0.96 12.22 2.12 ;
        RECT  10.86 1.52 12.22 1.68 ;
        RECT  11.02 1.84 11.30 2.12 ;
        RECT  11.02 0.96 11.30 1.24 ;
        RECT  11.02 0.96 11.18 2.12 ;
        RECT  10.86 1.46 11.18 1.74 ;
        END
    END QB
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.17  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.12 0.96 1.35 ;
        RECT  0.40 1.12 0.68 1.40 ;
        END
    END SEL
    PIN TD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.80 1.51 1.14 1.94 ;
        END
    END TD
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.06 1.46 2.40 1.80 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.78 1.33 4.06 1.70 ;
        END
    END CK
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 15.20 0.28 ;
        RECT  14.72 -0.28 15.02 0.32 ;
        RECT  14.66 0.64 14.94 0.92 ;
        RECT  14.72 -0.28 14.88 0.92 ;
        RECT  13.62 0.64 13.90 0.92 ;
        RECT  13.68 -0.28 13.84 0.92 ;
        RECT  12.58 0.64 12.86 0.92 ;
        RECT  12.64 -0.28 12.80 0.92 ;
        RECT  11.54 0.64 11.82 0.92 ;
        RECT  11.60 -0.28 11.76 0.92 ;
        RECT  10.50 0.64 10.78 0.92 ;
        RECT  10.56 -0.28 10.72 0.92 ;
        RECT  9.50 0.96 9.78 1.24 ;
        RECT  9.60 -0.28 9.76 1.24 ;
        RECT  6.78 0.68 7.06 0.96 ;
        RECT  6.84 -0.28 7.00 0.96 ;
        RECT  3.94 0.44 4.22 0.72 ;
        RECT  4.00 -0.28 4.16 0.72 ;
        RECT  2.30 0.68 2.58 0.96 ;
        RECT  2.36 -0.28 2.52 0.96 ;
        RECT  0.62 0.68 0.90 0.96 ;
        RECT  0.68 -0.28 0.84 0.96 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 15.20 3.48 ;
        RECT  14.72 2.88 15.02 3.48 ;
        RECT  14.66 2.16 14.94 2.44 ;
        RECT  14.72 2.16 14.88 3.48 ;
        RECT  13.62 2.16 13.90 2.44 ;
        RECT  13.68 2.16 13.84 3.48 ;
        RECT  12.58 2.16 12.86 2.44 ;
        RECT  12.64 2.16 12.80 3.48 ;
        RECT  11.54 2.16 11.82 2.44 ;
        RECT  11.60 2.16 11.76 3.48 ;
        RECT  10.50 2.03 10.78 2.31 ;
        RECT  10.56 2.03 10.72 3.48 ;
        RECT  9.50 2.62 9.78 3.48 ;
        RECT  6.78 1.92 7.06 2.20 ;
        RECT  6.84 1.92 7.00 3.48 ;
        RECT  3.90 2.62 4.18 3.48 ;
        RECT  2.30 2.04 2.58 2.32 ;
        RECT  2.36 2.04 2.52 3.48 ;
        RECT  0.60 2.62 0.88 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.08 0.68 0.38 0.96 ;
        RECT  0.08 0.68 0.24 2.32 ;
        RECT  0.08 2.04 0.38 2.32 ;
        RECT  0.08 2.16 1.28 2.32 ;
        RECT  1.12 2.16 1.28 2.64 ;
        RECT  1.28 2.48 1.56 2.76 ;
        RECT  1.46 0.68 1.74 0.96 ;
        RECT  1.52 1.12 2.88 1.28 ;
        RECT  2.60 1.12 2.88 1.40 ;
        RECT  1.52 0.68 1.68 2.32 ;
        RECT  1.46 2.04 1.74 2.32 ;
        RECT  3.40 0.44 3.70 0.72 ;
        RECT  3.40 0.94 4.40 1.10 ;
        RECT  4.12 0.88 4.40 1.16 ;
        RECT  3.40 0.44 3.56 2.14 ;
        RECT  3.40 1.86 3.70 2.14 ;
        RECT  4.46 0.44 4.74 0.72 ;
        RECT  4.58 1.40 4.88 1.68 ;
        RECT  4.58 0.44 4.74 2.14 ;
        RECT  4.46 1.86 4.74 2.14 ;
        RECT  2.82 0.68 3.20 0.96 ;
        RECT  4.94 0.68 5.22 0.96 ;
        RECT  5.04 0.68 5.20 2.20 ;
        RECT  3.04 0.68 3.20 2.46 ;
        RECT  4.94 1.92 5.22 2.20 ;
        RECT  4.94 1.92 5.10 2.46 ;
        RECT  2.82 2.04 3.20 2.32 ;
        RECT  3.04 2.30 5.10 2.46 ;
        RECT  5.46 0.68 5.74 0.96 ;
        RECT  5.46 1.92 5.74 2.20 ;
        RECT  5.52 0.68 5.68 2.70 ;
        RECT  6.12 2.42 6.40 2.70 ;
        RECT  5.52 2.54 6.40 2.70 ;
        RECT  6.12 0.68 6.40 0.96 ;
        RECT  6.18 0.68 6.34 2.20 ;
        RECT  6.12 1.92 6.40 2.20 ;
        RECT  7.30 0.68 7.58 0.96 ;
        RECT  6.64 1.44 7.52 1.60 ;
        RECT  6.64 1.38 6.92 1.66 ;
        RECT  7.36 0.68 7.52 2.20 ;
        RECT  7.30 1.92 7.58 2.20 ;
        RECT  7.98 0.44 9.44 0.60 ;
        RECT  9.16 0.44 9.44 0.80 ;
        RECT  7.98 0.44 8.14 1.04 ;
        RECT  7.86 0.76 8.14 1.04 ;
        RECT  7.88 0.76 8.04 2.20 ;
        RECT  7.82 1.92 8.10 2.20 ;
        RECT  8.98 0.96 9.26 1.24 ;
        RECT  8.98 1.46 9.98 1.62 ;
        RECT  9.70 1.40 9.98 1.68 ;
        RECT  8.98 0.96 9.14 2.12 ;
        RECT  8.98 1.84 9.26 2.12 ;
        RECT  8.38 0.76 8.66 1.04 ;
        RECT  10.02 0.96 10.30 1.24 ;
        RECT  10.02 1.84 10.30 2.12 ;
        RECT  8.40 0.76 8.56 2.20 ;
        RECT  8.34 1.92 8.62 2.20 ;
        RECT  8.46 1.92 8.62 2.44 ;
        RECT  10.14 0.96 10.30 2.72 ;
        RECT  8.46 2.28 10.30 2.44 ;
        RECT  10.12 2.44 10.40 2.72 ;
    END
END DFFDZSP8V1_0

MACRO DFFDZSP4V1_1
    CLASS CORE ;
    FOREIGN DFFDZSP4V1_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 21.15  LAYER ME1  ;
        ANTENNADIFFAREA 9.89  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.05  LAYER ME1  ;
        ANTENNAMAXAREACAR 20.22  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.97 1.46 10.34 1.74 ;
        RECT  9.85 1.84 10.13 2.12 ;
        RECT  9.97 0.96 10.13 2.12 ;
        RECT  9.85 0.96 10.13 1.24 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 21.15  LAYER ME1  ;
        ANTENNADIFFAREA 9.89  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.05  LAYER ME1  ;
        ANTENNAMAXAREACAR 20.22  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.89 1.84 11.17 2.12 ;
        RECT  10.89 0.96 11.17 1.24 ;
        RECT  10.89 0.96 11.14 2.12 ;
        RECT  10.86 1.46 11.14 1.74 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.24  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 18.44  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.81 1.19 2.25 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  0.91 0.81 1.19 1.09 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.86 1.46 3.37 1.74 ;
        END
    END CK
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END SEL
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.92  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 13.64  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.07 1.46 2.32 1.74 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.81 2.23 2.25 ;
        RECT  1.95 0.81 2.23 1.09 ;
        END
    END TD
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 12.00 3.48 ;
        RECT  11.47 2.88 11.82 3.48 ;
        RECT  11.41 2.16 11.69 2.44 ;
        RECT  11.47 2.16 11.63 3.48 ;
        RECT  10.37 2.16 10.65 2.44 ;
        RECT  10.43 2.16 10.59 3.48 ;
        RECT  9.33 1.84 9.61 2.12 ;
        RECT  9.39 1.84 9.55 3.48 ;
        RECT  8.33 2.62 8.61 3.48 ;
        RECT  5.77 1.92 6.05 2.20 ;
        RECT  5.83 1.92 5.99 3.48 ;
        RECT  2.95 2.62 3.23 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 12.00 0.28 ;
        RECT  11.47 -0.28 11.82 0.32 ;
        RECT  11.41 0.64 11.69 0.92 ;
        RECT  11.47 -0.28 11.63 0.92 ;
        RECT  10.37 0.64 10.65 0.92 ;
        RECT  10.43 -0.28 10.59 0.92 ;
        RECT  9.33 0.64 9.61 0.92 ;
        RECT  9.39 -0.28 9.55 0.92 ;
        RECT  8.33 0.96 8.61 1.24 ;
        RECT  8.43 -0.28 8.59 1.24 ;
        RECT  5.59 0.72 5.87 1.00 ;
        RECT  5.65 -0.28 5.81 1.00 ;
        RECT  2.95 0.87 3.23 1.15 ;
        RECT  3.01 -0.28 3.17 1.15 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  1.55 1.97 1.71 2.58 ;
        RECT  2.39 2.30 2.67 2.58 ;
        RECT  1.55 2.42 2.67 2.58 ;
        RECT  3.47 0.87 3.77 1.15 ;
        RECT  3.61 1.25 3.89 1.53 ;
        RECT  3.61 0.87 3.77 2.14 ;
        RECT  3.49 1.86 3.77 2.14 ;
        RECT  3.97 0.72 4.25 1.00 ;
        RECT  2.43 0.87 2.71 1.15 ;
        RECT  2.54 0.87 2.70 2.14 ;
        RECT  4.05 0.72 4.21 2.20 ;
        RECT  2.43 1.86 2.71 2.14 ;
        RECT  2.43 1.98 3.07 2.14 ;
        RECT  3.97 1.92 4.25 2.20 ;
        RECT  2.91 1.98 3.07 2.46 ;
        RECT  3.97 1.92 4.13 2.46 ;
        RECT  2.91 2.30 4.13 2.46 ;
        RECT  5.05 0.72 5.35 1.00 ;
        RECT  5.05 0.72 5.21 2.20 ;
        RECT  5.01 1.92 5.29 2.20 ;
        RECT  4.49 0.72 4.77 1.00 ;
        RECT  5.85 1.48 6.13 1.76 ;
        RECT  5.45 1.60 6.13 1.76 ;
        RECT  4.55 0.72 4.71 2.20 ;
        RECT  4.49 1.92 4.77 2.20 ;
        RECT  4.61 1.92 4.77 2.52 ;
        RECT  5.45 1.60 5.61 2.52 ;
        RECT  4.61 2.36 5.61 2.52 ;
        RECT  6.11 0.72 6.45 1.00 ;
        RECT  5.37 1.16 6.45 1.32 ;
        RECT  5.37 1.16 5.65 1.44 ;
        RECT  6.29 0.72 6.45 2.20 ;
        RECT  6.29 1.92 6.57 2.20 ;
        RECT  6.79 0.44 8.27 0.60 ;
        RECT  7.99 0.44 8.27 0.80 ;
        RECT  6.67 0.76 6.95 1.04 ;
        RECT  6.79 0.44 6.95 2.20 ;
        RECT  6.79 1.92 7.09 2.20 ;
        RECT  7.81 0.96 8.09 1.24 ;
        RECT  7.81 1.46 8.78 1.62 ;
        RECT  8.50 1.40 8.78 1.68 ;
        RECT  7.81 0.96 7.97 2.12 ;
        RECT  7.81 1.84 8.09 2.12 ;
        RECT  7.19 0.76 7.49 1.04 ;
        RECT  8.85 0.96 9.13 1.24 ;
        RECT  8.85 1.84 9.13 2.12 ;
        RECT  7.33 0.76 7.49 2.20 ;
        RECT  7.45 1.92 7.61 2.44 ;
        RECT  8.94 0.96 9.10 2.70 ;
        RECT  7.45 2.28 9.10 2.44 ;
        RECT  8.94 2.42 9.23 2.70 ;
    END
END DFFDZSP4V1_1

MACRO DFFDZSP4V1_0
    CLASS CORE ;
    FOREIGN DFFDZSP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 13.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.78 1.33 4.06 1.70 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.06 1.46 2.40 1.80 ;
        END
    END D
    PIN TD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.80 1.51 1.14 1.94 ;
        END
    END TD
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.17  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.12 0.96 1.35 ;
        RECT  0.40 1.12 0.68 1.40 ;
        END
    END SEL
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 23.99  LAYER ME1  ;
        ANTENNADIFFAREA 11.23  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.35  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.79  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.02 1.84 11.30 2.12 ;
        RECT  11.02 0.96 11.30 1.24 ;
        RECT  11.02 0.96 11.18 2.12 ;
        RECT  10.86 1.46 11.18 1.74 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 23.74  LAYER ME1  ;
        ANTENNADIFFAREA 11.23  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.35  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.60  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.06 1.84 12.34 2.12 ;
        RECT  12.06 0.96 12.34 1.24 ;
        RECT  12.12 0.96 12.28 2.12 ;
        END
    END Q
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 13.20 3.48 ;
        RECT  12.64 2.88 13.02 3.48 ;
        RECT  12.58 2.16 12.86 2.44 ;
        RECT  12.64 2.16 12.80 3.48 ;
        RECT  11.54 2.16 11.82 2.44 ;
        RECT  11.60 2.16 11.76 3.48 ;
        RECT  10.50 2.03 10.78 2.31 ;
        RECT  10.56 2.03 10.72 3.48 ;
        RECT  9.50 2.62 9.78 3.48 ;
        RECT  6.78 1.92 7.06 2.20 ;
        RECT  6.84 1.92 7.00 3.48 ;
        RECT  3.90 2.62 4.18 3.48 ;
        RECT  2.30 2.04 2.58 2.32 ;
        RECT  2.36 2.04 2.52 3.48 ;
        RECT  0.60 2.62 0.88 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 13.20 0.28 ;
        RECT  12.64 -0.28 13.02 0.32 ;
        RECT  12.58 0.64 12.86 0.92 ;
        RECT  12.64 -0.28 12.80 0.92 ;
        RECT  11.54 0.64 11.82 0.92 ;
        RECT  11.60 -0.28 11.76 0.92 ;
        RECT  10.50 0.64 10.78 0.92 ;
        RECT  10.56 -0.28 10.72 0.92 ;
        RECT  9.50 0.96 9.78 1.24 ;
        RECT  9.60 -0.28 9.76 1.24 ;
        RECT  6.78 0.68 7.06 0.96 ;
        RECT  6.84 -0.28 7.00 0.96 ;
        RECT  3.94 0.44 4.22 0.72 ;
        RECT  4.00 -0.28 4.16 0.72 ;
        RECT  2.30 0.68 2.58 0.96 ;
        RECT  2.36 -0.28 2.52 0.96 ;
        RECT  0.62 0.68 0.90 0.96 ;
        RECT  0.68 -0.28 0.84 0.96 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.08 0.68 0.38 0.96 ;
        RECT  0.08 0.68 0.24 2.32 ;
        RECT  0.08 2.04 0.38 2.32 ;
        RECT  0.08 2.16 1.28 2.32 ;
        RECT  1.12 2.16 1.28 2.64 ;
        RECT  1.28 2.48 1.56 2.76 ;
        RECT  1.46 0.68 1.74 0.96 ;
        RECT  1.52 1.12 2.88 1.28 ;
        RECT  2.60 1.12 2.88 1.40 ;
        RECT  1.52 0.68 1.68 2.32 ;
        RECT  1.46 2.04 1.74 2.32 ;
        RECT  3.40 0.44 3.70 0.72 ;
        RECT  3.40 0.94 4.40 1.10 ;
        RECT  4.12 0.88 4.40 1.16 ;
        RECT  3.40 0.44 3.56 2.14 ;
        RECT  3.40 1.86 3.70 2.14 ;
        RECT  4.46 0.44 4.74 0.72 ;
        RECT  4.58 1.40 4.88 1.68 ;
        RECT  4.58 0.44 4.74 2.14 ;
        RECT  4.46 1.86 4.74 2.14 ;
        RECT  2.82 0.68 3.20 0.96 ;
        RECT  4.94 0.68 5.22 0.96 ;
        RECT  5.04 0.68 5.20 2.20 ;
        RECT  3.04 0.68 3.20 2.46 ;
        RECT  4.94 1.92 5.22 2.20 ;
        RECT  4.94 1.92 5.10 2.46 ;
        RECT  2.82 2.04 3.20 2.32 ;
        RECT  3.04 2.30 5.10 2.46 ;
        RECT  5.46 0.68 5.74 0.96 ;
        RECT  5.46 1.92 5.74 2.20 ;
        RECT  5.52 0.68 5.68 2.70 ;
        RECT  6.12 2.42 6.40 2.70 ;
        RECT  5.52 2.54 6.40 2.70 ;
        RECT  6.12 0.68 6.40 0.96 ;
        RECT  6.18 0.68 6.34 2.20 ;
        RECT  6.12 1.92 6.40 2.20 ;
        RECT  7.30 0.68 7.58 0.96 ;
        RECT  6.64 1.44 7.52 1.60 ;
        RECT  6.64 1.38 6.92 1.66 ;
        RECT  7.36 0.68 7.52 2.20 ;
        RECT  7.30 1.92 7.58 2.20 ;
        RECT  7.98 0.44 9.44 0.60 ;
        RECT  9.16 0.44 9.44 0.80 ;
        RECT  7.98 0.44 8.14 1.04 ;
        RECT  7.86 0.76 8.14 1.04 ;
        RECT  7.88 0.76 8.04 2.20 ;
        RECT  7.82 1.92 8.10 2.20 ;
        RECT  8.98 0.96 9.26 1.24 ;
        RECT  8.98 1.46 9.98 1.62 ;
        RECT  9.70 1.40 9.98 1.68 ;
        RECT  8.98 0.96 9.14 2.12 ;
        RECT  8.98 1.84 9.26 2.12 ;
        RECT  8.38 0.76 8.66 1.04 ;
        RECT  10.02 0.96 10.30 1.24 ;
        RECT  10.02 1.84 10.30 2.12 ;
        RECT  8.40 0.76 8.56 2.20 ;
        RECT  8.34 1.92 8.62 2.20 ;
        RECT  8.46 1.92 8.62 2.44 ;
        RECT  10.14 0.96 10.30 2.72 ;
        RECT  8.46 2.28 10.30 2.44 ;
        RECT  10.12 2.44 10.40 2.72 ;
    END
END DFFDZSP4V1_0

MACRO DFFDZSP2V1_1
    CLASS CORE ;
    FOREIGN DFFDZSP2V1_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 18.90  LAYER ME1  ;
        ANTENNADIFFAREA 8.51  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.76  LAYER ME1  ;
        ANTENNAMAXAREACAR 24.92  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.33 1.84 9.61 2.12 ;
        RECT  9.33 0.96 9.61 1.24 ;
        RECT  9.33 0.96 9.54 2.12 ;
        RECT  9.26 1.46 9.54 1.74 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 19.20  LAYER ME1  ;
        ANTENNADIFFAREA 8.51  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.76  LAYER ME1  ;
        ANTENNAMAXAREACAR 25.32  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.37 1.84 10.65 2.12 ;
        RECT  10.37 0.96 10.65 1.24 ;
        RECT  10.37 0.96 10.53 2.12 ;
        RECT  10.06 1.46 10.53 1.74 ;
        END
    END Q
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.92  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 13.64  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.07 1.46 2.32 1.74 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.81 2.23 2.25 ;
        RECT  1.95 0.81 2.23 1.09 ;
        END
    END TD
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END SEL
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.86 1.46 3.37 1.74 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.24  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 18.44  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.81 1.19 2.25 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  0.91 0.81 1.19 1.09 ;
        END
    END D
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 10.80 0.28 ;
        RECT  10.34 -0.28 10.62 0.32 ;
        RECT  9.85 0.64 10.13 0.92 ;
        RECT  9.91 -0.28 10.07 0.92 ;
        RECT  8.33 0.96 8.61 1.24 ;
        RECT  8.43 -0.28 8.59 1.24 ;
        RECT  5.59 0.72 5.87 1.00 ;
        RECT  5.65 -0.28 5.81 1.00 ;
        RECT  2.95 0.87 3.23 1.15 ;
        RECT  3.01 -0.28 3.17 1.15 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 10.80 3.48 ;
        RECT  10.34 2.88 10.62 3.48 ;
        RECT  9.85 2.16 10.13 2.44 ;
        RECT  9.91 2.16 10.07 3.48 ;
        RECT  8.33 2.62 8.61 3.48 ;
        RECT  5.77 1.92 6.05 2.20 ;
        RECT  5.83 1.92 5.99 3.48 ;
        RECT  2.95 2.62 3.23 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  1.55 1.97 1.71 2.58 ;
        RECT  2.39 2.30 2.67 2.58 ;
        RECT  1.55 2.42 2.67 2.58 ;
        RECT  3.47 0.87 3.77 1.15 ;
        RECT  3.61 1.25 3.89 1.53 ;
        RECT  3.61 0.87 3.77 2.14 ;
        RECT  3.49 1.86 3.77 2.14 ;
        RECT  3.97 0.72 4.25 1.00 ;
        RECT  2.43 0.87 2.71 1.15 ;
        RECT  2.54 0.87 2.70 2.14 ;
        RECT  4.05 0.72 4.21 2.20 ;
        RECT  2.43 1.86 2.71 2.14 ;
        RECT  2.43 1.98 3.07 2.14 ;
        RECT  3.97 1.92 4.25 2.20 ;
        RECT  2.91 1.98 3.07 2.46 ;
        RECT  3.97 1.92 4.13 2.46 ;
        RECT  2.91 2.30 4.13 2.46 ;
        RECT  5.05 0.72 5.35 1.00 ;
        RECT  5.05 0.72 5.21 2.20 ;
        RECT  5.01 1.92 5.29 2.20 ;
        RECT  4.49 0.72 4.77 1.00 ;
        RECT  5.85 1.48 6.13 1.76 ;
        RECT  5.45 1.60 6.13 1.76 ;
        RECT  4.55 0.72 4.71 2.20 ;
        RECT  4.49 1.92 4.77 2.20 ;
        RECT  4.61 1.92 4.77 2.52 ;
        RECT  5.45 1.60 5.61 2.52 ;
        RECT  4.61 2.36 5.61 2.52 ;
        RECT  6.11 0.72 6.45 1.00 ;
        RECT  5.37 1.16 6.45 1.32 ;
        RECT  5.37 1.16 5.65 1.44 ;
        RECT  6.29 0.72 6.45 2.20 ;
        RECT  6.29 1.92 6.57 2.20 ;
        RECT  6.79 0.44 8.27 0.60 ;
        RECT  7.99 0.44 8.27 0.80 ;
        RECT  6.67 0.76 6.95 1.04 ;
        RECT  6.79 0.44 6.95 2.20 ;
        RECT  6.79 1.92 7.09 2.20 ;
        RECT  7.81 0.96 8.09 1.24 ;
        RECT  7.81 1.46 8.78 1.62 ;
        RECT  8.50 1.40 8.78 1.68 ;
        RECT  7.81 0.96 7.97 2.12 ;
        RECT  7.81 1.84 8.09 2.12 ;
        RECT  7.19 0.76 7.49 1.04 ;
        RECT  8.85 0.96 9.13 1.24 ;
        RECT  8.85 1.84 9.13 2.12 ;
        RECT  7.33 0.76 7.49 2.20 ;
        RECT  7.45 1.92 7.61 2.44 ;
        RECT  8.94 0.96 9.10 2.70 ;
        RECT  7.45 2.28 9.10 2.44 ;
        RECT  8.94 2.42 9.23 2.70 ;
    END
END DFFDZSP2V1_1

MACRO DFFDZSP2V1_0
    CLASS CORE ;
    FOREIGN DFFDZSP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 22.04  LAYER ME1  ;
        ANTENNADIFFAREA 9.88  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.06  LAYER ME1  ;
        ANTENNAMAXAREACAR 20.78  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.54 1.84 11.88 2.12 ;
        RECT  11.72 0.96 11.88 2.12 ;
        RECT  11.54 0.96 11.88 1.24 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 21.79  LAYER ME1  ;
        ANTENNADIFFAREA 9.88  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.06  LAYER ME1  ;
        ANTENNAMAXAREACAR 20.54  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.50 1.84 10.78 2.12 ;
        RECT  10.50 0.96 10.78 1.24 ;
        RECT  10.52 0.96 10.68 2.12 ;
        END
    END QB
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.17  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.12 0.96 1.35 ;
        RECT  0.40 1.12 0.68 1.40 ;
        END
    END SEL
    PIN TD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.80 1.51 1.14 1.94 ;
        END
    END TD
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.06 1.46 2.40 1.80 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.78 1.33 4.06 1.70 ;
        END
    END CK
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 12.00 0.28 ;
        RECT  11.54 -0.28 11.82 0.32 ;
        RECT  11.02 0.64 11.30 0.92 ;
        RECT  11.08 -0.28 11.24 0.92 ;
        RECT  9.50 0.96 9.78 1.24 ;
        RECT  9.60 -0.28 9.76 1.24 ;
        RECT  6.78 0.68 7.06 0.96 ;
        RECT  6.84 -0.28 7.00 0.96 ;
        RECT  3.94 0.44 4.22 0.72 ;
        RECT  4.00 -0.28 4.16 0.72 ;
        RECT  2.30 0.68 2.58 0.96 ;
        RECT  2.36 -0.28 2.52 0.96 ;
        RECT  0.62 0.68 0.90 0.96 ;
        RECT  0.68 -0.28 0.84 0.96 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 12.00 3.48 ;
        RECT  11.54 2.88 11.82 3.48 ;
        RECT  11.02 2.16 11.30 2.44 ;
        RECT  11.08 2.16 11.24 3.48 ;
        RECT  9.50 2.62 9.78 3.48 ;
        RECT  6.78 1.92 7.06 2.20 ;
        RECT  6.84 1.92 7.00 3.48 ;
        RECT  3.90 2.62 4.18 3.48 ;
        RECT  2.30 2.04 2.58 2.32 ;
        RECT  2.36 2.04 2.52 3.48 ;
        RECT  0.60 2.62 0.88 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.08 0.68 0.38 0.96 ;
        RECT  0.08 0.68 0.24 2.32 ;
        RECT  0.08 2.04 0.38 2.32 ;
        RECT  0.08 2.16 1.28 2.32 ;
        RECT  1.12 2.16 1.28 2.64 ;
        RECT  1.28 2.48 1.56 2.76 ;
        RECT  1.46 0.68 1.74 0.96 ;
        RECT  1.52 1.12 2.88 1.28 ;
        RECT  2.60 1.12 2.88 1.40 ;
        RECT  1.52 0.68 1.68 2.32 ;
        RECT  1.46 2.04 1.74 2.32 ;
        RECT  3.40 0.44 3.70 0.72 ;
        RECT  3.40 0.94 4.40 1.10 ;
        RECT  4.12 0.88 4.40 1.16 ;
        RECT  3.40 0.44 3.56 2.14 ;
        RECT  3.40 1.86 3.70 2.14 ;
        RECT  4.46 0.44 4.74 0.72 ;
        RECT  4.58 1.40 4.88 1.68 ;
        RECT  4.58 0.44 4.74 2.14 ;
        RECT  4.46 1.86 4.74 2.14 ;
        RECT  2.82 0.68 3.20 0.96 ;
        RECT  4.94 0.68 5.22 0.96 ;
        RECT  5.04 0.68 5.20 2.20 ;
        RECT  3.04 0.68 3.20 2.46 ;
        RECT  4.94 1.92 5.22 2.20 ;
        RECT  4.94 1.92 5.10 2.46 ;
        RECT  2.82 2.04 3.20 2.32 ;
        RECT  3.04 2.30 5.10 2.46 ;
        RECT  5.46 0.68 5.74 0.96 ;
        RECT  5.46 1.92 5.74 2.20 ;
        RECT  5.52 0.68 5.68 2.70 ;
        RECT  6.12 2.42 6.40 2.70 ;
        RECT  5.52 2.54 6.40 2.70 ;
        RECT  6.12 0.68 6.40 0.96 ;
        RECT  6.18 0.68 6.34 2.20 ;
        RECT  6.12 1.92 6.40 2.20 ;
        RECT  7.30 0.68 7.58 0.96 ;
        RECT  6.64 1.44 7.52 1.60 ;
        RECT  6.64 1.38 6.92 1.66 ;
        RECT  7.36 0.68 7.52 2.20 ;
        RECT  7.30 1.92 7.58 2.20 ;
        RECT  7.98 0.44 9.44 0.60 ;
        RECT  9.16 0.44 9.44 0.80 ;
        RECT  7.98 0.44 8.14 1.04 ;
        RECT  7.86 0.76 8.14 1.04 ;
        RECT  7.88 0.76 8.04 2.20 ;
        RECT  7.82 1.92 8.10 2.20 ;
        RECT  8.98 0.96 9.26 1.24 ;
        RECT  8.98 1.46 9.98 1.62 ;
        RECT  9.70 1.40 9.98 1.68 ;
        RECT  8.98 0.96 9.14 2.12 ;
        RECT  8.98 1.84 9.26 2.12 ;
        RECT  8.38 0.76 8.66 1.04 ;
        RECT  10.02 0.96 10.30 1.24 ;
        RECT  10.02 1.84 10.30 2.12 ;
        RECT  8.40 0.76 8.56 2.20 ;
        RECT  8.34 1.92 8.62 2.20 ;
        RECT  8.46 1.92 8.62 2.44 ;
        RECT  10.14 0.96 10.30 2.72 ;
        RECT  8.46 2.28 10.30 2.44 ;
        RECT  10.12 2.44 10.40 2.72 ;
    END
END DFFDZSP2V1_0

MACRO DFFDZSP1V1_1
    CLASS CORE ;
    FOREIGN DFFDZSP1V1_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.24  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 18.44  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.81 1.19 2.25 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  0.91 0.81 1.19 1.09 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.87 1.46 3.37 1.74 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 18.99  LAYER ME1  ;
        ANTENNADIFFAREA 7.82  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.60  LAYER ME1  ;
        ANTENNAMAXAREACAR 31.41  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.33 1.90 9.61 2.18 ;
        RECT  9.33 0.96 9.61 1.24 ;
        RECT  9.33 0.96 9.49 2.18 ;
        RECT  9.26 1.46 9.49 1.74 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 19.28  LAYER ME1  ;
        ANTENNADIFFAREA 7.82  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.60  LAYER ME1  ;
        ANTENNAMAXAREACAR 31.87  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.37 1.90 10.65 2.18 ;
        RECT  10.37 0.96 10.65 1.24 ;
        RECT  10.37 0.96 10.53 2.18 ;
        RECT  10.06 1.46 10.53 1.74 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END SEL
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.92  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 13.64  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.07 1.46 2.32 1.74 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.81 2.23 2.25 ;
        RECT  1.95 0.81 2.23 1.09 ;
        END
    END TD
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 10.80 3.48 ;
        RECT  10.34 2.88 10.62 3.48 ;
        RECT  9.85 1.90 10.13 2.18 ;
        RECT  9.91 1.90 10.07 3.48 ;
        RECT  8.33 2.62 8.61 3.48 ;
        RECT  5.77 1.92 6.05 2.20 ;
        RECT  5.83 1.92 5.99 3.48 ;
        RECT  2.95 2.62 3.23 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 10.80 0.28 ;
        RECT  10.34 -0.28 10.62 0.32 ;
        RECT  9.85 0.96 10.13 1.24 ;
        RECT  9.91 -0.28 10.07 1.24 ;
        RECT  8.33 0.96 8.61 1.24 ;
        RECT  8.43 -0.28 8.59 1.24 ;
        RECT  5.59 0.72 5.87 1.00 ;
        RECT  5.65 -0.28 5.81 1.00 ;
        RECT  2.95 0.87 3.23 1.15 ;
        RECT  3.01 -0.28 3.17 1.15 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  1.55 1.97 1.71 2.58 ;
        RECT  2.39 2.30 2.67 2.58 ;
        RECT  1.55 2.42 2.67 2.58 ;
        RECT  3.47 0.87 3.77 1.15 ;
        RECT  3.61 1.25 3.89 1.53 ;
        RECT  3.61 0.87 3.77 2.14 ;
        RECT  3.49 1.86 3.77 2.14 ;
        RECT  3.97 0.72 4.25 1.00 ;
        RECT  2.43 0.87 2.71 1.15 ;
        RECT  4.05 0.72 4.21 2.20 ;
        RECT  2.55 0.87 2.71 2.14 ;
        RECT  2.43 1.86 2.71 2.14 ;
        RECT  2.43 1.98 3.07 2.14 ;
        RECT  3.97 1.92 4.25 2.20 ;
        RECT  2.91 1.98 3.07 2.46 ;
        RECT  3.97 1.92 4.13 2.46 ;
        RECT  2.91 2.30 4.13 2.46 ;
        RECT  5.05 0.72 5.35 1.00 ;
        RECT  5.05 0.72 5.21 2.20 ;
        RECT  5.01 1.92 5.29 2.20 ;
        RECT  4.49 0.72 4.77 1.00 ;
        RECT  5.85 1.48 6.13 1.76 ;
        RECT  5.45 1.60 6.13 1.76 ;
        RECT  4.55 0.72 4.71 2.20 ;
        RECT  4.49 1.92 4.77 2.20 ;
        RECT  4.61 1.92 4.77 2.52 ;
        RECT  5.45 1.60 5.61 2.52 ;
        RECT  4.61 2.36 5.61 2.52 ;
        RECT  6.11 0.72 6.45 1.00 ;
        RECT  5.37 1.16 6.45 1.32 ;
        RECT  5.37 1.16 5.65 1.44 ;
        RECT  6.29 0.72 6.45 2.20 ;
        RECT  6.29 1.92 6.57 2.20 ;
        RECT  6.79 0.44 8.27 0.60 ;
        RECT  7.99 0.44 8.27 0.80 ;
        RECT  6.67 0.76 6.95 1.04 ;
        RECT  6.79 0.44 6.95 2.20 ;
        RECT  6.79 1.92 7.09 2.20 ;
        RECT  7.81 0.96 8.09 1.24 ;
        RECT  7.81 1.46 8.75 1.62 ;
        RECT  8.47 1.40 8.75 1.68 ;
        RECT  7.81 0.96 7.97 2.12 ;
        RECT  7.81 1.84 8.09 2.12 ;
        RECT  7.19 0.76 7.49 1.04 ;
        RECT  8.85 0.96 9.13 1.24 ;
        RECT  8.85 1.84 9.13 2.12 ;
        RECT  7.33 0.76 7.49 2.20 ;
        RECT  7.45 1.92 7.61 2.44 ;
        RECT  8.94 0.96 9.10 2.70 ;
        RECT  7.45 2.28 9.10 2.44 ;
        RECT  8.94 2.42 9.23 2.70 ;
    END
END DFFDZSP1V1_1

MACRO DFFDZSP1V1_0
    CLASS CORE ;
    FOREIGN DFFDZSP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 21.90  LAYER ME1  ;
        ANTENNADIFFAREA 9.19  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.91  LAYER ME1  ;
        ANTENNAMAXAREACAR 24.14  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.50 1.84 10.78 2.12 ;
        RECT  10.50 0.96 10.78 1.24 ;
        RECT  10.52 0.96 10.68 2.12 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 22.15  LAYER ME1  ;
        ANTENNADIFFAREA 9.19  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.91  LAYER ME1  ;
        ANTENNAMAXAREACAR 24.42  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.54 1.84 11.88 2.12 ;
        RECT  11.72 0.96 11.88 2.12 ;
        RECT  11.54 0.96 11.88 1.24 ;
        END
    END Q
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.78 1.33 4.06 1.70 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.06 1.46 2.40 1.80 ;
        END
    END D
    PIN TD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.80 1.51 1.14 1.94 ;
        END
    END TD
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.17  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.12 0.96 1.35 ;
        RECT  0.40 1.12 0.68 1.40 ;
        END
    END SEL
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 12.00 3.48 ;
        RECT  11.54 2.88 11.82 3.48 ;
        RECT  11.02 1.84 11.30 2.12 ;
        RECT  11.08 1.84 11.24 3.48 ;
        RECT  9.50 2.62 9.78 3.48 ;
        RECT  6.78 1.92 7.06 2.20 ;
        RECT  6.84 1.92 7.00 3.48 ;
        RECT  3.90 2.62 4.18 3.48 ;
        RECT  2.30 2.04 2.58 2.32 ;
        RECT  2.36 2.04 2.52 3.48 ;
        RECT  0.60 2.62 0.88 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 12.00 0.28 ;
        RECT  11.54 -0.28 11.82 0.32 ;
        RECT  11.02 0.96 11.30 1.24 ;
        RECT  11.08 -0.28 11.24 1.24 ;
        RECT  9.50 0.96 9.78 1.24 ;
        RECT  9.60 -0.28 9.76 1.24 ;
        RECT  6.78 0.68 7.06 0.96 ;
        RECT  6.84 -0.28 7.00 0.96 ;
        RECT  3.94 0.44 4.22 0.72 ;
        RECT  4.00 -0.28 4.16 0.72 ;
        RECT  2.30 0.68 2.58 0.96 ;
        RECT  2.36 -0.28 2.52 0.96 ;
        RECT  0.62 0.68 0.90 0.96 ;
        RECT  0.68 -0.28 0.84 0.96 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.08 0.68 0.38 0.96 ;
        RECT  0.08 0.68 0.24 2.32 ;
        RECT  0.08 2.04 0.38 2.32 ;
        RECT  0.08 2.16 1.28 2.32 ;
        RECT  1.12 2.16 1.28 2.64 ;
        RECT  1.28 2.48 1.56 2.76 ;
        RECT  1.46 0.68 1.74 0.96 ;
        RECT  1.52 1.12 2.88 1.28 ;
        RECT  2.60 1.12 2.88 1.40 ;
        RECT  1.52 0.68 1.68 2.32 ;
        RECT  1.46 2.04 1.74 2.32 ;
        RECT  3.40 0.44 3.70 0.72 ;
        RECT  3.40 0.94 4.40 1.10 ;
        RECT  4.12 0.88 4.40 1.16 ;
        RECT  3.40 0.44 3.56 2.14 ;
        RECT  3.40 1.86 3.70 2.14 ;
        RECT  4.46 0.44 4.74 0.72 ;
        RECT  4.58 1.40 4.88 1.68 ;
        RECT  4.58 0.44 4.74 2.14 ;
        RECT  4.46 1.86 4.74 2.14 ;
        RECT  2.82 0.68 3.20 0.96 ;
        RECT  4.94 0.68 5.22 0.96 ;
        RECT  5.04 0.68 5.20 2.20 ;
        RECT  3.04 0.68 3.20 2.46 ;
        RECT  4.94 1.92 5.22 2.20 ;
        RECT  4.94 1.92 5.10 2.46 ;
        RECT  2.82 2.04 3.20 2.32 ;
        RECT  3.04 2.30 5.10 2.46 ;
        RECT  5.46 0.68 5.74 0.96 ;
        RECT  5.46 1.92 5.74 2.20 ;
        RECT  5.52 0.68 5.68 2.70 ;
        RECT  6.12 2.42 6.40 2.70 ;
        RECT  5.52 2.54 6.40 2.70 ;
        RECT  6.12 0.68 6.40 0.96 ;
        RECT  6.18 0.68 6.34 2.20 ;
        RECT  6.12 1.92 6.40 2.20 ;
        RECT  7.30 0.68 7.58 0.96 ;
        RECT  6.64 1.44 7.52 1.60 ;
        RECT  6.64 1.38 6.92 1.66 ;
        RECT  7.36 0.68 7.52 2.20 ;
        RECT  7.30 1.92 7.58 2.20 ;
        RECT  7.98 0.44 9.44 0.60 ;
        RECT  9.16 0.44 9.44 0.80 ;
        RECT  7.98 0.44 8.14 1.04 ;
        RECT  7.86 0.76 8.14 1.04 ;
        RECT  7.88 0.76 8.04 2.20 ;
        RECT  7.82 1.92 8.10 2.20 ;
        RECT  8.98 0.96 9.26 1.24 ;
        RECT  8.98 1.46 9.98 1.62 ;
        RECT  9.70 1.40 9.98 1.68 ;
        RECT  8.98 0.96 9.14 2.12 ;
        RECT  8.98 1.84 9.26 2.12 ;
        RECT  8.38 0.76 8.66 1.04 ;
        RECT  10.02 0.96 10.30 1.24 ;
        RECT  10.02 1.84 10.30 2.12 ;
        RECT  8.40 0.76 8.56 2.20 ;
        RECT  8.34 1.92 8.62 2.20 ;
        RECT  8.46 1.92 8.62 2.44 ;
        RECT  10.14 0.96 10.30 2.44 ;
        RECT  8.46 2.28 10.54 2.44 ;
        RECT  10.26 2.28 10.54 2.62 ;
    END
END DFFDZSP1V1_0

MACRO DFFDSZSP8V1_0
    CLASS CORE ;
    FOREIGN DFFDSZSP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 31.16  LAYER ME1  ;
        ANTENNADIFFAREA 14.98  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.62  LAYER ME1  ;
        ANTENNAMAXAREACAR 19.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  15.25 1.90 15.53 2.50 ;
        RECT  15.25 0.64 15.53 1.24 ;
        RECT  15.25 0.64 15.41 2.50 ;
        RECT  14.33 1.52 15.41 1.68 ;
        RECT  14.33 1.46 14.74 1.74 ;
        RECT  14.21 1.90 14.49 2.50 ;
        RECT  14.33 0.64 14.49 2.50 ;
        RECT  14.21 0.64 14.49 1.24 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 31.16  LAYER ME1  ;
        ANTENNADIFFAREA 14.95  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.62  LAYER ME1  ;
        ANTENNAMAXAREACAR 19.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.17 1.90 13.45 2.50 ;
        RECT  13.17 0.64 13.45 1.24 ;
        RECT  13.17 0.64 13.33 2.50 ;
        RECT  12.06 1.52 13.33 1.68 ;
        RECT  12.13 1.90 12.41 2.50 ;
        RECT  12.13 0.64 12.41 1.24 ;
        RECT  12.13 0.64 12.34 2.50 ;
        RECT  12.06 1.46 12.34 1.74 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.20  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.83  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.81 1.19 2.25 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  0.91 0.81 1.19 1.09 ;
        END
    END D
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END SEL
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.87  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 12.90  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.06 1.46 2.34 1.74 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.81 2.23 2.25 ;
        RECT  1.95 0.81 2.23 1.09 ;
        END
    END TD
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.53 1.40 9.95 1.68 ;
        END
    END SB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.24 1.40 3.54 1.76 ;
        END
    END CK
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 16.40 0.28 ;
        RECT  15.83 -0.28 16.22 0.32 ;
        RECT  15.77 0.64 16.05 1.24 ;
        RECT  15.83 -0.28 15.99 1.24 ;
        RECT  14.73 0.64 15.01 1.24 ;
        RECT  14.79 -0.28 14.95 1.24 ;
        RECT  13.69 0.64 13.97 1.24 ;
        RECT  13.75 -0.28 13.91 1.24 ;
        RECT  12.65 0.64 12.93 1.24 ;
        RECT  12.71 -0.28 12.87 1.24 ;
        RECT  11.61 0.64 11.89 1.24 ;
        RECT  11.67 -0.28 11.83 1.24 ;
        RECT  10.61 0.88 10.89 1.16 ;
        RECT  10.67 -0.28 10.83 1.16 ;
        RECT  9.13 -0.28 9.41 0.68 ;
        RECT  2.71 -0.28 2.99 0.68 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 16.40 3.48 ;
        RECT  15.83 2.88 16.22 3.48 ;
        RECT  15.77 1.90 16.05 2.50 ;
        RECT  15.83 1.90 15.99 3.48 ;
        RECT  14.73 1.90 15.01 2.50 ;
        RECT  14.79 1.90 14.95 3.48 ;
        RECT  13.69 1.90 13.97 2.50 ;
        RECT  13.75 1.90 13.91 3.48 ;
        RECT  12.65 1.90 12.93 2.50 ;
        RECT  12.71 1.90 12.87 3.48 ;
        RECT  11.61 1.90 11.89 2.50 ;
        RECT  11.67 1.90 11.83 3.48 ;
        RECT  10.37 2.40 10.65 3.48 ;
        RECT  9.57 1.84 9.85 2.12 ;
        RECT  9.63 1.84 9.79 3.48 ;
        RECT  8.57 1.84 8.85 2.12 ;
        RECT  8.63 1.84 8.79 3.48 ;
        RECT  7.57 1.84 7.85 2.12 ;
        RECT  7.67 1.84 7.83 3.48 ;
        RECT  2.71 2.52 2.99 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  1.55 1.97 1.71 2.57 ;
        RECT  1.55 2.41 2.37 2.57 ;
        RECT  2.09 2.41 2.37 2.69 ;
        RECT  3.47 0.96 3.86 1.24 ;
        RECT  3.70 1.46 4.02 1.74 ;
        RECT  3.70 0.95 3.86 2.19 ;
        RECT  3.47 1.92 3.75 2.20 ;
        RECT  4.07 0.44 4.35 0.72 ;
        RECT  3.15 0.56 4.35 0.72 ;
        RECT  3.15 0.56 3.31 1.12 ;
        RECT  2.43 0.96 3.31 1.12 ;
        RECT  2.43 0.96 2.71 1.24 ;
        RECT  2.55 0.96 2.71 2.20 ;
        RECT  2.43 1.92 2.71 2.20 ;
        RECT  2.43 2.04 3.31 2.20 ;
        RECT  3.15 2.04 3.31 2.64 ;
        RECT  3.15 2.48 4.25 2.64 ;
        RECT  3.97 2.48 4.25 2.76 ;
        RECT  5.59 0.76 5.91 1.04 ;
        RECT  5.59 0.76 5.75 2.00 ;
        RECT  5.25 1.84 6.29 2.00 ;
        RECT  5.25 1.84 5.53 2.12 ;
        RECT  6.01 1.84 6.29 2.12 ;
        RECT  6.15 0.76 6.43 1.04 ;
        RECT  6.27 0.76 6.43 1.36 ;
        RECT  7.11 1.08 7.39 1.36 ;
        RECT  6.27 1.20 7.39 1.36 ;
        RECT  6.53 1.20 6.69 2.12 ;
        RECT  6.53 1.84 6.81 2.12 ;
        RECT  4.63 0.86 4.91 1.14 ;
        RECT  4.07 0.98 4.91 1.14 ;
        RECT  4.07 0.96 4.35 1.24 ;
        RECT  4.29 0.98 4.45 2.12 ;
        RECT  4.41 1.84 4.57 2.44 ;
        RECT  4.41 2.28 7.51 2.44 ;
        RECT  7.23 2.28 7.51 2.56 ;
        RECT  6.67 0.76 7.95 0.92 ;
        RECT  6.67 0.76 6.95 1.04 ;
        RECT  7.67 0.76 7.95 1.16 ;
        RECT  7.67 0.76 7.83 1.68 ;
        RECT  8.71 1.40 8.99 1.68 ;
        RECT  7.25 1.52 8.99 1.68 ;
        RECT  8.01 1.52 8.17 2.12 ;
        RECT  7.25 1.52 7.41 2.12 ;
        RECT  7.05 1.84 7.41 2.12 ;
        RECT  8.01 1.84 8.37 2.12 ;
        RECT  5.27 0.44 8.87 0.60 ;
        RECT  8.71 0.44 8.87 1.04 ;
        RECT  8.71 0.88 9.37 1.04 ;
        RECT  5.27 0.44 5.43 1.14 ;
        RECT  9.09 0.88 9.37 1.16 ;
        RECT  5.15 0.86 5.31 1.46 ;
        RECT  4.93 1.30 5.31 1.46 ;
        RECT  9.15 0.88 9.31 2.12 ;
        RECT  4.93 1.30 5.09 2.12 ;
        RECT  4.81 1.84 5.09 2.12 ;
        RECT  9.09 1.84 9.37 2.12 ;
        RECT  9.71 0.88 9.99 1.16 ;
        RECT  9.71 1.00 10.27 1.16 ;
        RECT  10.11 1.00 10.27 2.12 ;
        RECT  10.09 1.84 10.37 2.12 ;
        RECT  10.09 1.96 10.97 2.12 ;
        RECT  10.81 1.96 10.97 2.64 ;
        RECT  10.81 2.48 11.44 2.64 ;
        RECT  11.16 2.48 11.44 2.76 ;
        RECT  11.13 0.88 11.41 1.16 ;
        RECT  10.43 1.46 11.55 1.62 ;
        RECT  10.43 1.40 10.71 1.68 ;
        RECT  11.25 1.40 11.55 1.68 ;
        RECT  11.25 0.88 11.41 2.12 ;
        RECT  11.13 1.84 11.41 2.12 ;
    END
END DFFDSZSP8V1_0

MACRO DFFDSZSP4V1_0
    CLASS CORE ;
    FOREIGN DFFDSZSP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.24 1.40 3.54 1.76 ;
        END
    END CK
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.53 1.40 9.95 1.68 ;
        END
    END SB
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.87  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 12.90  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.06 1.46 2.34 1.74 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.81 2.23 2.25 ;
        RECT  1.95 0.81 2.23 1.09 ;
        END
    END TD
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END SEL
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.20  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.83  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.81 1.19 2.25 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  0.91 0.81 1.19 1.09 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 26.88  LAYER ME1  ;
        ANTENNADIFFAREA 11.91  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.05  LAYER ME1  ;
        ANTENNAMAXAREACAR 25.68  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.13 1.90 12.41 2.50 ;
        RECT  12.13 0.64 12.41 1.24 ;
        RECT  12.13 0.64 12.34 2.50 ;
        RECT  12.06 1.46 12.34 1.74 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 26.88  LAYER ME1  ;
        ANTENNADIFFAREA 11.94  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.05  LAYER ME1  ;
        ANTENNAMAXAREACAR 25.68  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.26 1.46 13.54 1.74 ;
        RECT  13.17 1.90 13.45 2.50 ;
        RECT  13.26 0.64 13.45 2.50 ;
        RECT  13.17 0.64 13.45 1.24 ;
        END
    END QB
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 14.40 3.48 ;
        RECT  13.78 2.88 14.22 3.48 ;
        RECT  13.69 1.90 13.97 2.50 ;
        RECT  13.78 1.90 13.94 3.48 ;
        RECT  12.65 1.90 12.93 2.50 ;
        RECT  12.71 1.90 12.87 3.48 ;
        RECT  11.61 1.90 11.89 2.50 ;
        RECT  11.67 1.90 11.83 3.48 ;
        RECT  10.37 2.40 10.65 3.48 ;
        RECT  9.57 1.84 9.85 2.12 ;
        RECT  9.63 1.84 9.79 3.48 ;
        RECT  8.57 1.84 8.85 2.12 ;
        RECT  8.63 1.84 8.79 3.48 ;
        RECT  7.57 1.84 7.85 2.12 ;
        RECT  7.67 1.84 7.83 3.48 ;
        RECT  2.71 2.52 2.99 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 14.40 0.28 ;
        RECT  13.78 -0.28 14.22 0.32 ;
        RECT  13.69 0.64 13.97 1.24 ;
        RECT  13.78 -0.28 13.94 1.24 ;
        RECT  12.65 0.64 12.93 1.24 ;
        RECT  12.71 -0.28 12.87 1.24 ;
        RECT  11.61 0.64 11.89 1.24 ;
        RECT  11.67 -0.28 11.83 1.24 ;
        RECT  10.61 0.88 10.89 1.16 ;
        RECT  10.67 -0.28 10.83 1.16 ;
        RECT  9.13 -0.28 9.41 0.68 ;
        RECT  2.71 -0.28 2.99 0.68 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  1.55 1.97 1.71 2.57 ;
        RECT  1.55 2.41 2.37 2.57 ;
        RECT  2.09 2.41 2.37 2.69 ;
        RECT  3.47 0.96 3.86 1.24 ;
        RECT  3.70 1.46 4.02 1.74 ;
        RECT  3.70 0.95 3.86 2.19 ;
        RECT  3.47 1.92 3.75 2.20 ;
        RECT  4.07 0.44 4.35 0.72 ;
        RECT  3.15 0.56 4.35 0.72 ;
        RECT  3.15 0.56 3.31 1.12 ;
        RECT  2.43 0.96 3.31 1.12 ;
        RECT  2.43 0.96 2.71 1.24 ;
        RECT  2.55 0.96 2.71 2.20 ;
        RECT  2.43 1.92 2.71 2.20 ;
        RECT  2.43 2.04 3.31 2.20 ;
        RECT  3.15 2.04 3.31 2.64 ;
        RECT  3.15 2.48 4.25 2.64 ;
        RECT  3.97 2.48 4.25 2.76 ;
        RECT  5.59 0.76 5.91 1.04 ;
        RECT  5.59 0.76 5.75 2.00 ;
        RECT  5.25 1.84 6.29 2.00 ;
        RECT  5.25 1.84 5.53 2.12 ;
        RECT  6.01 1.84 6.29 2.12 ;
        RECT  6.15 0.76 6.43 1.04 ;
        RECT  6.27 0.76 6.43 1.36 ;
        RECT  7.11 1.08 7.39 1.36 ;
        RECT  6.27 1.20 7.39 1.36 ;
        RECT  6.53 1.20 6.69 2.12 ;
        RECT  6.53 1.84 6.81 2.12 ;
        RECT  4.63 0.86 4.91 1.14 ;
        RECT  4.07 0.98 4.91 1.14 ;
        RECT  4.07 0.96 4.35 1.24 ;
        RECT  4.29 0.98 4.45 2.12 ;
        RECT  4.41 1.84 4.57 2.44 ;
        RECT  4.41 2.28 7.51 2.44 ;
        RECT  7.23 2.28 7.51 2.56 ;
        RECT  6.67 0.76 7.95 0.92 ;
        RECT  6.67 0.76 6.95 1.04 ;
        RECT  7.67 0.76 7.95 1.16 ;
        RECT  7.67 0.76 7.83 1.68 ;
        RECT  8.71 1.40 8.99 1.68 ;
        RECT  7.25 1.52 8.99 1.68 ;
        RECT  8.01 1.52 8.17 2.12 ;
        RECT  7.25 1.52 7.41 2.12 ;
        RECT  7.05 1.84 7.41 2.12 ;
        RECT  8.01 1.84 8.37 2.12 ;
        RECT  5.27 0.44 8.87 0.60 ;
        RECT  8.71 0.44 8.87 1.04 ;
        RECT  8.71 0.88 9.37 1.04 ;
        RECT  5.27 0.44 5.43 1.14 ;
        RECT  9.09 0.88 9.37 1.16 ;
        RECT  5.15 0.86 5.31 1.46 ;
        RECT  4.93 1.30 5.31 1.46 ;
        RECT  9.15 0.88 9.31 2.12 ;
        RECT  4.93 1.30 5.09 2.12 ;
        RECT  4.81 1.84 5.09 2.12 ;
        RECT  9.09 1.84 9.37 2.12 ;
        RECT  9.71 0.88 9.99 1.16 ;
        RECT  9.71 1.00 10.27 1.16 ;
        RECT  10.11 1.00 10.27 2.12 ;
        RECT  10.09 1.84 10.37 2.12 ;
        RECT  10.09 1.96 10.97 2.12 ;
        RECT  10.81 1.96 10.97 2.64 ;
        RECT  10.81 2.48 11.44 2.64 ;
        RECT  11.16 2.48 11.44 2.76 ;
        RECT  11.13 0.88 11.41 1.16 ;
        RECT  10.43 1.46 11.55 1.62 ;
        RECT  10.43 1.40 10.71 1.68 ;
        RECT  11.25 1.40 11.55 1.68 ;
        RECT  11.25 0.88 11.41 2.12 ;
        RECT  11.13 1.84 11.41 2.12 ;
    END
END DFFDSZSP4V1_0

MACRO DFFDSZSP2V1_0
    CLASS CORE ;
    FOREIGN DFFDSZSP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 13.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 24.69  LAYER ME1  ;
        ANTENNADIFFAREA 10.36  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.76  LAYER ME1  ;
        ANTENNAMAXAREACAR 32.56  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.77 1.46 13.12 1.74 ;
        RECT  12.65 1.90 12.93 2.50 ;
        RECT  12.77 0.64 12.93 2.50 ;
        RECT  12.65 0.64 12.93 1.24 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 24.69  LAYER ME1  ;
        ANTENNADIFFAREA 10.36  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.76  LAYER ME1  ;
        ANTENNAMAXAREACAR 32.56  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.73 1.46 12.34 1.74 ;
        RECT  11.61 1.90 11.89 2.50 ;
        RECT  11.73 0.64 11.89 2.50 ;
        RECT  11.61 0.64 11.89 1.24 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.20  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.83  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.81 1.19 2.25 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  0.91 0.81 1.19 1.09 ;
        END
    END D
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END SEL
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.87  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 12.90  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.06 1.46 2.34 1.74 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.81 2.23 2.25 ;
        RECT  1.95 0.81 2.23 1.09 ;
        END
    END TD
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.53 1.40 9.95 1.68 ;
        END
    END SB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.24 1.40 3.54 1.76 ;
        END
    END CK
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 13.20 0.28 ;
        RECT  12.74 -0.28 13.02 0.32 ;
        RECT  12.13 0.64 12.41 1.24 ;
        RECT  12.19 -0.28 12.35 1.24 ;
        RECT  10.61 0.88 10.89 1.16 ;
        RECT  10.67 -0.28 10.83 1.16 ;
        RECT  9.13 -0.28 9.41 0.68 ;
        RECT  2.71 -0.28 2.99 0.68 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 13.20 3.48 ;
        RECT  12.74 2.88 13.02 3.48 ;
        RECT  12.13 1.90 12.41 2.50 ;
        RECT  12.19 1.90 12.35 3.48 ;
        RECT  10.37 2.40 10.65 3.48 ;
        RECT  9.57 1.84 9.85 2.12 ;
        RECT  9.63 1.84 9.79 3.48 ;
        RECT  8.57 1.84 8.85 2.12 ;
        RECT  8.63 1.84 8.79 3.48 ;
        RECT  7.57 1.84 7.85 2.12 ;
        RECT  7.67 1.84 7.83 3.48 ;
        RECT  2.71 2.52 2.99 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  1.55 1.97 1.71 2.57 ;
        RECT  1.55 2.41 2.37 2.57 ;
        RECT  2.09 2.41 2.37 2.69 ;
        RECT  3.47 0.96 3.86 1.24 ;
        RECT  3.70 1.46 4.02 1.74 ;
        RECT  3.70 0.95 3.86 2.19 ;
        RECT  3.47 1.92 3.75 2.20 ;
        RECT  4.07 0.44 4.35 0.72 ;
        RECT  3.15 0.56 4.35 0.72 ;
        RECT  3.15 0.56 3.31 1.12 ;
        RECT  2.43 0.96 3.31 1.12 ;
        RECT  2.43 0.96 2.71 1.24 ;
        RECT  2.55 0.96 2.71 2.20 ;
        RECT  2.43 1.92 2.71 2.20 ;
        RECT  2.43 2.04 3.31 2.20 ;
        RECT  3.15 2.04 3.31 2.64 ;
        RECT  3.15 2.48 4.25 2.64 ;
        RECT  3.97 2.48 4.25 2.76 ;
        RECT  5.59 0.76 5.91 1.04 ;
        RECT  5.59 0.76 5.75 2.00 ;
        RECT  5.25 1.84 6.29 2.00 ;
        RECT  5.25 1.84 5.53 2.12 ;
        RECT  6.01 1.84 6.29 2.12 ;
        RECT  6.15 0.76 6.43 1.04 ;
        RECT  6.27 0.76 6.43 1.36 ;
        RECT  7.11 1.08 7.39 1.36 ;
        RECT  6.27 1.20 7.39 1.36 ;
        RECT  6.53 1.20 6.69 2.12 ;
        RECT  6.53 1.84 6.81 2.12 ;
        RECT  4.63 0.86 4.91 1.14 ;
        RECT  4.07 0.98 4.91 1.14 ;
        RECT  4.07 0.96 4.35 1.24 ;
        RECT  4.29 0.98 4.45 2.12 ;
        RECT  4.41 1.84 4.57 2.44 ;
        RECT  4.41 2.28 7.51 2.44 ;
        RECT  7.23 2.28 7.51 2.56 ;
        RECT  6.67 0.76 7.95 0.92 ;
        RECT  6.67 0.76 6.95 1.04 ;
        RECT  7.67 0.76 7.95 1.16 ;
        RECT  7.67 0.76 7.83 1.68 ;
        RECT  8.71 1.40 8.99 1.68 ;
        RECT  7.25 1.52 8.99 1.68 ;
        RECT  8.01 1.52 8.17 2.12 ;
        RECT  7.25 1.52 7.41 2.12 ;
        RECT  7.05 1.84 7.41 2.12 ;
        RECT  8.01 1.84 8.37 2.12 ;
        RECT  5.27 0.44 8.87 0.60 ;
        RECT  8.71 0.44 8.87 1.04 ;
        RECT  8.71 0.88 9.37 1.04 ;
        RECT  5.27 0.44 5.43 1.14 ;
        RECT  9.09 0.88 9.37 1.16 ;
        RECT  5.15 0.86 5.31 1.46 ;
        RECT  4.93 1.30 5.31 1.46 ;
        RECT  9.15 0.88 9.31 2.12 ;
        RECT  4.93 1.30 5.09 2.12 ;
        RECT  4.81 1.84 5.09 2.12 ;
        RECT  9.09 1.84 9.37 2.12 ;
        RECT  9.71 0.88 9.99 1.16 ;
        RECT  9.71 1.00 10.27 1.16 ;
        RECT  10.11 1.00 10.27 2.12 ;
        RECT  10.09 1.84 10.37 2.12 ;
        RECT  10.09 1.96 10.97 2.12 ;
        RECT  10.81 1.96 10.97 2.64 ;
        RECT  10.81 2.48 11.44 2.64 ;
        RECT  11.16 2.48 11.44 2.76 ;
        RECT  11.13 0.88 11.41 1.16 ;
        RECT  10.43 1.46 11.55 1.62 ;
        RECT  10.43 1.40 10.71 1.68 ;
        RECT  11.25 1.40 11.55 1.68 ;
        RECT  11.25 0.88 11.41 2.12 ;
        RECT  11.13 1.84 11.41 2.12 ;
    END
END DFFDSZSP2V1_0

MACRO DFFDSZSP1V1_0
    CLASS CORE ;
    FOREIGN DFFDSZSP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 13.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.20  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.83  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.81 1.19 2.25 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  0.91 0.81 1.19 1.09 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.24 1.40 3.54 1.76 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 23.94  LAYER ME1  ;
        ANTENNADIFFAREA 9.67  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.60  LAYER ME1  ;
        ANTENNAMAXAREACAR 39.59  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.77 1.46 13.12 1.74 ;
        RECT  12.65 1.90 12.93 2.18 ;
        RECT  12.77 0.96 12.93 2.18 ;
        RECT  12.65 0.96 12.93 1.24 ;
        END
    END QB
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.53 1.40 9.95 1.68 ;
        END
    END SB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 24.26  LAYER ME1  ;
        ANTENNADIFFAREA 9.67  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.60  LAYER ME1  ;
        ANTENNAMAXAREACAR 40.11  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.73 1.46 12.34 1.74 ;
        RECT  11.61 1.90 11.89 2.18 ;
        RECT  11.73 0.96 11.89 2.18 ;
        RECT  11.61 0.96 11.89 1.24 ;
        END
    END Q
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.87  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 12.90  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.06 1.46 2.34 1.74 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.81 2.23 2.25 ;
        RECT  1.95 0.81 2.23 1.09 ;
        END
    END TD
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END SEL
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 13.20 0.28 ;
        RECT  12.74 -0.28 13.02 0.32 ;
        RECT  12.13 0.96 12.41 1.24 ;
        RECT  12.19 -0.28 12.35 1.24 ;
        RECT  10.61 0.88 10.89 1.16 ;
        RECT  10.67 -0.28 10.83 1.16 ;
        RECT  9.13 -0.28 9.41 0.68 ;
        RECT  2.71 -0.28 2.99 0.68 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 13.20 3.48 ;
        RECT  12.74 2.88 13.02 3.48 ;
        RECT  12.13 1.90 12.41 2.18 ;
        RECT  12.19 1.90 12.35 3.48 ;
        RECT  10.37 2.40 10.65 3.48 ;
        RECT  9.57 1.84 9.85 2.12 ;
        RECT  9.63 1.84 9.79 3.48 ;
        RECT  8.57 1.84 8.85 2.12 ;
        RECT  8.63 1.84 8.79 3.48 ;
        RECT  7.57 1.84 7.85 2.12 ;
        RECT  7.67 1.84 7.83 3.48 ;
        RECT  2.71 2.52 2.99 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  1.55 1.97 1.71 2.57 ;
        RECT  1.55 2.41 2.37 2.57 ;
        RECT  2.09 2.41 2.37 2.69 ;
        RECT  3.47 0.96 3.86 1.24 ;
        RECT  3.70 1.46 4.02 1.74 ;
        RECT  3.70 0.95 3.86 2.19 ;
        RECT  3.47 1.92 3.75 2.20 ;
        RECT  4.07 0.44 4.35 0.72 ;
        RECT  3.15 0.56 4.35 0.72 ;
        RECT  3.15 0.56 3.31 1.12 ;
        RECT  2.43 0.96 3.31 1.12 ;
        RECT  2.43 0.96 2.71 1.24 ;
        RECT  2.55 0.96 2.71 2.20 ;
        RECT  2.43 1.92 2.71 2.20 ;
        RECT  2.43 2.04 3.31 2.20 ;
        RECT  3.15 2.04 3.31 2.64 ;
        RECT  3.15 2.48 4.25 2.64 ;
        RECT  3.97 2.48 4.25 2.76 ;
        RECT  5.59 0.76 5.91 1.04 ;
        RECT  5.59 0.76 5.75 2.00 ;
        RECT  5.25 1.84 6.29 2.00 ;
        RECT  5.25 1.84 5.53 2.12 ;
        RECT  6.01 1.84 6.29 2.12 ;
        RECT  6.15 0.76 6.43 1.04 ;
        RECT  6.27 0.76 6.43 1.36 ;
        RECT  7.11 1.08 7.39 1.36 ;
        RECT  6.27 1.20 7.39 1.36 ;
        RECT  6.53 1.20 6.69 2.12 ;
        RECT  6.53 1.84 6.81 2.12 ;
        RECT  4.63 0.86 4.91 1.14 ;
        RECT  4.07 0.98 4.91 1.14 ;
        RECT  4.07 0.96 4.35 1.24 ;
        RECT  4.29 0.98 4.45 2.12 ;
        RECT  4.41 1.84 4.57 2.44 ;
        RECT  4.41 2.28 7.51 2.44 ;
        RECT  7.23 2.28 7.51 2.56 ;
        RECT  6.67 0.76 7.95 0.92 ;
        RECT  6.67 0.76 6.95 1.04 ;
        RECT  7.67 0.76 7.95 1.16 ;
        RECT  7.67 0.76 7.83 1.68 ;
        RECT  8.71 1.40 8.99 1.68 ;
        RECT  7.25 1.52 8.99 1.68 ;
        RECT  8.01 1.52 8.17 2.12 ;
        RECT  7.25 1.52 7.41 2.12 ;
        RECT  7.05 1.84 7.41 2.12 ;
        RECT  8.01 1.84 8.37 2.12 ;
        RECT  5.27 0.44 8.87 0.60 ;
        RECT  8.71 0.44 8.87 1.04 ;
        RECT  8.71 0.88 9.37 1.04 ;
        RECT  5.27 0.44 5.43 1.14 ;
        RECT  9.09 0.88 9.37 1.16 ;
        RECT  5.15 0.86 5.31 1.46 ;
        RECT  4.93 1.30 5.31 1.46 ;
        RECT  9.15 0.88 9.31 2.12 ;
        RECT  4.93 1.30 5.09 2.12 ;
        RECT  4.81 1.84 5.09 2.12 ;
        RECT  9.09 1.84 9.37 2.12 ;
        RECT  9.71 0.88 9.99 1.16 ;
        RECT  9.71 1.00 10.27 1.16 ;
        RECT  10.11 1.00 10.27 2.12 ;
        RECT  10.09 1.84 10.37 2.12 ;
        RECT  10.09 1.96 10.97 2.12 ;
        RECT  10.81 1.96 10.97 2.64 ;
        RECT  10.81 2.48 11.44 2.64 ;
        RECT  11.16 2.48 11.44 2.76 ;
        RECT  11.13 0.88 11.41 1.16 ;
        RECT  10.43 1.46 11.55 1.62 ;
        RECT  10.43 1.40 10.71 1.68 ;
        RECT  11.25 1.40 11.55 1.68 ;
        RECT  11.25 0.88 11.41 2.12 ;
        RECT  11.13 1.84 11.41 2.12 ;
    END
END DFFDSZSP1V1_0

MACRO DFFDSSP8V1_0
    CLASS CORE ;
    FOREIGN DFFDSSP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 27.83  LAYER ME1  ;
        ANTENNADIFFAREA 13.83  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.56  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.89  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.92 1.90 13.20 2.50 ;
        RECT  12.92 0.64 13.20 1.24 ;
        RECT  12.92 0.64 13.08 2.50 ;
        RECT  12.00 1.52 13.08 1.68 ;
        RECT  12.00 1.46 12.34 1.74 ;
        RECT  11.88 1.90 12.16 2.50 ;
        RECT  12.00 0.64 12.16 2.50 ;
        RECT  11.88 0.64 12.16 1.24 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 27.83  LAYER ME1  ;
        ANTENNADIFFAREA 13.80  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.56  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.89  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.84 1.90 11.12 2.50 ;
        RECT  10.84 0.64 11.12 1.24 ;
        RECT  10.84 0.64 11.00 2.50 ;
        RECT  9.92 1.52 11.00 1.68 ;
        RECT  9.92 1.46 10.34 1.74 ;
        RECT  9.80 1.90 10.08 2.50 ;
        RECT  9.92 0.64 10.08 2.50 ;
        RECT  9.80 0.64 10.08 1.24 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.18 1.40 7.60 1.68 ;
        END
    END SB
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.40 0.70 1.76 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.40 1.16 1.76 ;
        END
    END CK
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 14.00 0.28 ;
        RECT  13.50 -0.28 13.82 0.32 ;
        RECT  13.44 0.64 13.72 1.24 ;
        RECT  13.50 -0.28 13.66 1.24 ;
        RECT  12.40 0.64 12.68 1.24 ;
        RECT  12.46 -0.28 12.62 1.24 ;
        RECT  11.36 0.64 11.64 1.24 ;
        RECT  11.42 -0.28 11.58 1.24 ;
        RECT  10.32 0.64 10.60 1.24 ;
        RECT  10.38 -0.28 10.54 1.24 ;
        RECT  9.28 0.64 9.56 1.24 ;
        RECT  9.34 -0.28 9.50 1.24 ;
        RECT  8.28 0.88 8.56 1.16 ;
        RECT  8.34 -0.28 8.50 1.16 ;
        RECT  6.80 -0.28 7.08 0.68 ;
        RECT  0.38 -0.28 0.66 0.68 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 14.00 3.48 ;
        RECT  13.50 2.88 13.82 3.48 ;
        RECT  13.44 1.90 13.72 2.50 ;
        RECT  13.50 1.90 13.66 3.48 ;
        RECT  12.40 1.90 12.68 2.50 ;
        RECT  12.46 1.90 12.62 3.48 ;
        RECT  11.36 1.90 11.64 2.50 ;
        RECT  11.42 1.90 11.58 3.48 ;
        RECT  10.32 1.90 10.60 2.50 ;
        RECT  10.38 1.90 10.54 3.48 ;
        RECT  9.28 1.90 9.56 2.50 ;
        RECT  9.34 1.90 9.50 3.48 ;
        RECT  8.04 2.40 8.32 3.48 ;
        RECT  7.24 1.84 7.52 2.12 ;
        RECT  7.30 1.84 7.46 3.48 ;
        RECT  6.24 1.84 6.52 2.12 ;
        RECT  6.30 1.84 6.46 3.48 ;
        RECT  5.24 1.84 5.52 2.12 ;
        RECT  5.34 1.84 5.50 3.48 ;
        RECT  0.38 2.48 0.66 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  1.14 0.96 1.48 1.24 ;
        RECT  1.32 1.46 1.64 1.74 ;
        RECT  1.32 0.96 1.48 2.20 ;
        RECT  1.14 1.92 1.48 2.20 ;
        RECT  1.74 0.44 2.02 0.72 ;
        RECT  0.82 0.56 2.02 0.72 ;
        RECT  0.82 0.56 0.98 1.12 ;
        RECT  0.08 0.96 0.98 1.12 ;
        RECT  0.08 0.96 0.38 1.24 ;
        RECT  0.08 0.96 0.24 2.20 ;
        RECT  0.08 1.92 0.38 2.20 ;
        RECT  0.08 2.04 0.98 2.20 ;
        RECT  0.82 2.04 0.98 2.64 ;
        RECT  0.82 2.48 1.92 2.64 ;
        RECT  1.64 2.48 1.92 2.76 ;
        RECT  3.26 0.76 3.58 1.04 ;
        RECT  3.26 0.76 3.42 2.00 ;
        RECT  2.92 1.84 3.96 2.00 ;
        RECT  2.92 1.84 3.20 2.12 ;
        RECT  3.68 1.84 3.96 2.12 ;
        RECT  3.82 0.76 4.10 1.04 ;
        RECT  3.94 0.76 4.10 1.36 ;
        RECT  4.78 1.08 5.06 1.36 ;
        RECT  3.94 1.20 5.06 1.36 ;
        RECT  4.20 1.20 4.36 2.12 ;
        RECT  4.20 1.84 4.48 2.12 ;
        RECT  2.30 0.86 2.58 1.14 ;
        RECT  1.74 0.98 2.58 1.14 ;
        RECT  1.74 0.96 2.02 1.24 ;
        RECT  1.96 0.98 2.12 2.12 ;
        RECT  2.08 1.84 2.24 2.44 ;
        RECT  2.08 2.28 5.18 2.44 ;
        RECT  4.90 2.28 5.18 2.56 ;
        RECT  4.34 0.76 5.62 0.92 ;
        RECT  4.34 0.76 4.62 1.04 ;
        RECT  5.34 0.76 5.62 1.16 ;
        RECT  5.34 0.76 5.50 1.68 ;
        RECT  6.38 1.40 6.66 1.68 ;
        RECT  4.92 1.52 6.66 1.68 ;
        RECT  5.68 1.52 5.84 2.12 ;
        RECT  4.92 1.52 5.08 2.12 ;
        RECT  4.72 1.84 5.08 2.12 ;
        RECT  5.68 1.84 6.04 2.12 ;
        RECT  2.94 0.44 6.54 0.60 ;
        RECT  6.38 0.44 6.54 1.04 ;
        RECT  6.38 0.88 7.04 1.04 ;
        RECT  2.94 0.44 3.10 1.14 ;
        RECT  6.76 0.88 7.04 1.16 ;
        RECT  2.82 0.86 2.98 1.46 ;
        RECT  2.60 1.30 2.98 1.46 ;
        RECT  6.82 0.88 6.98 2.12 ;
        RECT  2.60 1.30 2.76 2.12 ;
        RECT  2.48 1.84 2.76 2.12 ;
        RECT  6.76 1.84 7.04 2.12 ;
        RECT  7.38 0.88 7.66 1.16 ;
        RECT  7.38 1.00 7.92 1.16 ;
        RECT  7.76 1.00 7.92 2.12 ;
        RECT  7.76 1.84 8.04 2.12 ;
        RECT  7.76 1.96 8.64 2.12 ;
        RECT  8.48 1.96 8.64 2.64 ;
        RECT  8.48 2.48 9.11 2.64 ;
        RECT  8.83 2.48 9.11 2.76 ;
        RECT  8.80 0.88 9.08 1.16 ;
        RECT  8.10 1.46 9.22 1.62 ;
        RECT  8.10 1.40 8.38 1.68 ;
        RECT  8.92 1.40 9.22 1.68 ;
        RECT  8.92 0.88 9.08 2.12 ;
        RECT  8.80 1.84 9.08 2.12 ;
    END
END DFFDSSP8V1_0

MACRO DFFDSSP4V1_0
    CLASS CORE ;
    FOREIGN DFFDSSP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.40 1.16 1.76 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.40 0.70 1.76 ;
        END
    END D
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.18 1.40 7.60 1.68 ;
        END
    END SB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 23.64  LAYER ME1  ;
        ANTENNADIFFAREA 10.76  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.98  LAYER ME1  ;
        ANTENNAMAXAREACAR 24.15  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.92 1.46 10.34 1.74 ;
        RECT  9.80 1.90 10.08 2.50 ;
        RECT  9.92 0.64 10.08 2.50 ;
        RECT  9.80 0.64 10.08 1.24 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 23.64  LAYER ME1  ;
        ANTENNADIFFAREA 10.79  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.98  LAYER ME1  ;
        ANTENNAMAXAREACAR 24.15  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.85 1.46 11.14 1.74 ;
        RECT  10.84 1.90 11.12 2.50 ;
        RECT  10.85 0.64 11.12 2.50 ;
        RECT  10.84 0.64 11.12 1.24 ;
        END
    END QB
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 12.00 3.48 ;
        RECT  11.42 2.88 11.82 3.48 ;
        RECT  11.36 1.90 11.64 2.50 ;
        RECT  11.42 1.90 11.58 3.48 ;
        RECT  10.32 1.90 10.60 2.50 ;
        RECT  10.38 1.90 10.54 3.48 ;
        RECT  9.28 1.90 9.56 2.50 ;
        RECT  9.34 1.90 9.50 3.48 ;
        RECT  8.04 2.40 8.32 3.48 ;
        RECT  7.24 1.84 7.52 2.12 ;
        RECT  7.30 1.84 7.46 3.48 ;
        RECT  6.24 1.84 6.52 2.12 ;
        RECT  6.30 1.84 6.46 3.48 ;
        RECT  5.24 1.84 5.52 2.12 ;
        RECT  5.34 1.84 5.50 3.48 ;
        RECT  0.38 2.48 0.66 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 12.00 0.28 ;
        RECT  11.42 -0.28 11.82 0.32 ;
        RECT  11.36 0.64 11.64 1.24 ;
        RECT  11.42 -0.28 11.58 1.24 ;
        RECT  10.32 0.64 10.60 1.24 ;
        RECT  10.38 -0.28 10.54 1.24 ;
        RECT  9.28 0.64 9.56 1.24 ;
        RECT  9.34 -0.28 9.50 1.24 ;
        RECT  8.28 0.88 8.56 1.16 ;
        RECT  8.34 -0.28 8.50 1.16 ;
        RECT  6.80 -0.28 7.08 0.68 ;
        RECT  0.38 -0.28 0.66 0.68 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  1.14 0.96 1.48 1.24 ;
        RECT  1.32 1.46 1.64 1.74 ;
        RECT  1.32 0.96 1.48 2.20 ;
        RECT  1.14 1.92 1.48 2.20 ;
        RECT  1.74 0.44 2.02 0.72 ;
        RECT  0.82 0.56 2.02 0.72 ;
        RECT  0.82 0.56 0.98 1.12 ;
        RECT  0.08 0.96 0.98 1.12 ;
        RECT  0.08 0.96 0.38 1.24 ;
        RECT  0.08 0.96 0.24 2.20 ;
        RECT  0.08 1.92 0.38 2.20 ;
        RECT  0.08 2.04 0.98 2.20 ;
        RECT  0.82 2.04 0.98 2.64 ;
        RECT  0.82 2.48 1.92 2.64 ;
        RECT  1.64 2.48 1.92 2.76 ;
        RECT  3.26 0.76 3.58 1.04 ;
        RECT  3.26 0.76 3.42 2.00 ;
        RECT  2.92 1.84 3.96 2.00 ;
        RECT  2.92 1.84 3.20 2.12 ;
        RECT  3.68 1.84 3.96 2.12 ;
        RECT  3.82 0.76 4.10 1.04 ;
        RECT  3.94 0.76 4.10 1.36 ;
        RECT  4.78 1.08 5.06 1.36 ;
        RECT  3.94 1.20 5.06 1.36 ;
        RECT  4.20 1.20 4.36 2.12 ;
        RECT  4.20 1.84 4.48 2.12 ;
        RECT  2.30 0.86 2.58 1.14 ;
        RECT  1.74 0.98 2.58 1.14 ;
        RECT  1.74 0.96 2.02 1.24 ;
        RECT  1.96 0.98 2.12 2.12 ;
        RECT  2.08 1.84 2.24 2.44 ;
        RECT  2.08 2.28 5.18 2.44 ;
        RECT  4.90 2.28 5.18 2.56 ;
        RECT  4.34 0.76 5.62 0.92 ;
        RECT  4.34 0.76 4.62 1.04 ;
        RECT  5.34 0.76 5.62 1.16 ;
        RECT  5.34 0.76 5.50 1.68 ;
        RECT  6.38 1.40 6.66 1.68 ;
        RECT  4.92 1.52 6.66 1.68 ;
        RECT  5.68 1.52 5.84 2.12 ;
        RECT  4.92 1.52 5.08 2.12 ;
        RECT  4.72 1.84 5.08 2.12 ;
        RECT  5.68 1.84 6.04 2.12 ;
        RECT  2.94 0.44 6.54 0.60 ;
        RECT  6.38 0.44 6.54 1.04 ;
        RECT  6.38 0.88 7.04 1.04 ;
        RECT  2.94 0.44 3.10 1.14 ;
        RECT  6.76 0.88 7.04 1.16 ;
        RECT  2.82 0.86 2.98 1.46 ;
        RECT  2.60 1.30 2.98 1.46 ;
        RECT  6.82 0.88 6.98 2.12 ;
        RECT  2.60 1.30 2.76 2.12 ;
        RECT  2.48 1.84 2.76 2.12 ;
        RECT  6.76 1.84 7.04 2.12 ;
        RECT  7.38 0.88 7.66 1.16 ;
        RECT  7.38 1.00 7.92 1.16 ;
        RECT  7.76 1.00 7.92 2.12 ;
        RECT  7.76 1.84 8.04 2.12 ;
        RECT  7.76 1.96 8.64 2.12 ;
        RECT  8.48 1.96 8.64 2.64 ;
        RECT  8.48 2.48 9.11 2.64 ;
        RECT  8.83 2.48 9.11 2.76 ;
        RECT  8.80 0.88 9.08 1.16 ;
        RECT  8.10 1.46 9.22 1.62 ;
        RECT  8.10 1.40 8.38 1.68 ;
        RECT  8.92 1.40 9.22 1.68 ;
        RECT  8.92 0.88 9.08 2.12 ;
        RECT  8.80 1.84 9.08 2.12 ;
    END
END DFFDSSP4V1_0

MACRO DFFDSSP2V1_0
    CLASS CORE ;
    FOREIGN DFFDSSP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 21.37  LAYER ME1  ;
        ANTENNADIFFAREA 9.21  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.69  LAYER ME1  ;
        ANTENNAMAXAREACAR 30.92  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.44 1.46 10.72 1.74 ;
        RECT  10.32 1.90 10.60 2.50 ;
        RECT  10.44 0.64 10.60 2.50 ;
        RECT  10.32 0.64 10.60 1.24 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 21.37  LAYER ME1  ;
        ANTENNADIFFAREA 9.21  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.69  LAYER ME1  ;
        ANTENNAMAXAREACAR 30.92  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.40 1.46 9.94 1.74 ;
        RECT  9.28 1.90 9.56 2.50 ;
        RECT  9.40 0.64 9.56 2.50 ;
        RECT  9.28 0.64 9.56 1.24 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.18 1.40 7.60 1.68 ;
        END
    END SB
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.40 0.70 1.76 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.40 1.16 1.76 ;
        END
    END CK
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 10.80 0.28 ;
        RECT  10.34 -0.28 10.62 0.32 ;
        RECT  9.80 0.64 10.08 1.24 ;
        RECT  9.86 -0.28 10.02 1.24 ;
        RECT  8.28 0.88 8.56 1.16 ;
        RECT  8.34 -0.28 8.50 1.16 ;
        RECT  6.80 -0.28 7.08 0.68 ;
        RECT  0.38 -0.28 0.66 0.68 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 10.80 3.48 ;
        RECT  10.34 2.88 10.62 3.48 ;
        RECT  9.80 1.90 10.08 2.50 ;
        RECT  9.86 1.90 10.02 3.48 ;
        RECT  8.04 2.40 8.32 3.48 ;
        RECT  7.24 1.84 7.52 2.12 ;
        RECT  7.30 1.84 7.46 3.48 ;
        RECT  6.24 1.84 6.52 2.12 ;
        RECT  6.30 1.84 6.46 3.48 ;
        RECT  5.24 1.84 5.52 2.12 ;
        RECT  5.34 1.84 5.50 3.48 ;
        RECT  0.38 2.48 0.66 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  1.14 0.96 1.48 1.24 ;
        RECT  1.32 1.46 1.64 1.74 ;
        RECT  1.32 0.96 1.48 2.20 ;
        RECT  1.14 1.92 1.48 2.20 ;
        RECT  1.74 0.44 2.02 0.72 ;
        RECT  0.82 0.56 2.02 0.72 ;
        RECT  0.82 0.56 0.98 1.12 ;
        RECT  0.08 0.96 0.98 1.12 ;
        RECT  0.08 0.96 0.38 1.24 ;
        RECT  0.08 0.96 0.24 2.20 ;
        RECT  0.08 1.92 0.38 2.20 ;
        RECT  0.08 2.04 0.98 2.20 ;
        RECT  0.82 2.04 0.98 2.64 ;
        RECT  0.82 2.48 1.92 2.64 ;
        RECT  1.64 2.48 1.92 2.76 ;
        RECT  3.26 0.76 3.58 1.04 ;
        RECT  3.26 0.76 3.42 2.00 ;
        RECT  2.92 1.84 3.96 2.00 ;
        RECT  2.92 1.84 3.20 2.12 ;
        RECT  3.68 1.84 3.96 2.12 ;
        RECT  3.82 0.76 4.10 1.04 ;
        RECT  3.94 0.76 4.10 1.36 ;
        RECT  4.78 1.08 5.06 1.36 ;
        RECT  3.94 1.20 5.06 1.36 ;
        RECT  4.20 1.20 4.36 2.12 ;
        RECT  4.20 1.84 4.48 2.12 ;
        RECT  2.30 0.86 2.58 1.14 ;
        RECT  1.74 0.98 2.58 1.14 ;
        RECT  1.74 0.96 2.02 1.24 ;
        RECT  1.96 0.98 2.12 2.12 ;
        RECT  2.08 1.84 2.24 2.44 ;
        RECT  2.08 2.28 5.18 2.44 ;
        RECT  4.90 2.28 5.18 2.56 ;
        RECT  4.34 0.76 5.62 0.92 ;
        RECT  4.34 0.76 4.62 1.04 ;
        RECT  5.34 0.76 5.62 1.16 ;
        RECT  5.34 0.76 5.50 1.68 ;
        RECT  6.38 1.40 6.66 1.68 ;
        RECT  4.92 1.52 6.66 1.68 ;
        RECT  5.68 1.52 5.84 2.12 ;
        RECT  4.92 1.52 5.08 2.12 ;
        RECT  4.72 1.84 5.08 2.12 ;
        RECT  5.68 1.84 6.04 2.12 ;
        RECT  2.94 0.44 6.54 0.60 ;
        RECT  6.38 0.44 6.54 1.04 ;
        RECT  6.38 0.88 7.04 1.04 ;
        RECT  2.94 0.44 3.10 1.14 ;
        RECT  6.76 0.88 7.04 1.16 ;
        RECT  2.82 0.86 2.98 1.46 ;
        RECT  2.60 1.30 2.98 1.46 ;
        RECT  6.82 0.88 6.98 2.12 ;
        RECT  2.60 1.30 2.76 2.12 ;
        RECT  2.48 1.84 2.76 2.12 ;
        RECT  6.76 1.84 7.04 2.12 ;
        RECT  7.38 0.88 7.66 1.16 ;
        RECT  7.38 1.00 7.92 1.16 ;
        RECT  7.76 1.00 7.92 2.12 ;
        RECT  7.76 1.84 8.04 2.12 ;
        RECT  7.76 1.96 8.64 2.12 ;
        RECT  8.48 1.96 8.64 2.64 ;
        RECT  8.48 2.48 9.11 2.64 ;
        RECT  8.83 2.48 9.11 2.76 ;
        RECT  8.80 0.88 9.08 1.16 ;
        RECT  8.10 1.46 9.22 1.62 ;
        RECT  8.10 1.40 8.38 1.68 ;
        RECT  8.92 1.40 9.22 1.68 ;
        RECT  8.92 0.88 9.08 2.12 ;
        RECT  8.80 1.84 9.08 2.12 ;
    END
END DFFDSSP2V1_0

MACRO DFFDSSP1V1_0
    CLASS CORE ;
    FOREIGN DFFDSSP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 20.64  LAYER ME1  ;
        ANTENNADIFFAREA 8.51  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.54  LAYER ME1  ;
        ANTENNAMAXAREACAR 38.39  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.44 1.46 10.72 1.74 ;
        RECT  10.32 1.90 10.60 2.18 ;
        RECT  10.44 0.96 10.60 2.18 ;
        RECT  10.32 0.96 10.60 1.24 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 20.93  LAYER ME1  ;
        ANTENNADIFFAREA 8.51  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.54  LAYER ME1  ;
        ANTENNAMAXAREACAR 38.94  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.40 1.46 9.94 1.74 ;
        RECT  9.28 1.90 9.56 2.18 ;
        RECT  9.40 0.96 9.56 2.18 ;
        RECT  9.28 0.96 9.56 1.24 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.40 0.70 1.76 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.40 1.16 1.76 ;
        END
    END CK
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.18 1.40 7.60 1.68 ;
        END
    END SB
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 10.80 3.48 ;
        RECT  10.34 2.88 10.62 3.48 ;
        RECT  9.80 1.90 10.08 2.18 ;
        RECT  9.86 1.90 10.02 3.48 ;
        RECT  8.04 2.40 8.32 3.48 ;
        RECT  7.24 1.84 7.52 2.12 ;
        RECT  7.30 1.84 7.46 3.48 ;
        RECT  6.24 1.84 6.52 2.12 ;
        RECT  6.30 1.84 6.46 3.48 ;
        RECT  5.24 1.84 5.52 2.12 ;
        RECT  5.34 1.84 5.50 3.48 ;
        RECT  0.38 2.48 0.66 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 10.80 0.28 ;
        RECT  10.34 -0.28 10.62 0.32 ;
        RECT  9.80 0.96 10.08 1.24 ;
        RECT  9.86 -0.28 10.02 1.24 ;
        RECT  8.28 0.88 8.56 1.16 ;
        RECT  8.34 -0.28 8.50 1.16 ;
        RECT  6.80 -0.28 7.08 0.68 ;
        RECT  0.38 -0.28 0.66 0.68 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  1.14 0.96 1.48 1.24 ;
        RECT  1.32 1.46 1.64 1.74 ;
        RECT  1.32 0.96 1.48 2.20 ;
        RECT  1.14 1.92 1.48 2.20 ;
        RECT  1.74 0.44 2.02 0.72 ;
        RECT  0.82 0.56 2.02 0.72 ;
        RECT  0.82 0.56 0.98 1.12 ;
        RECT  0.08 0.96 0.98 1.12 ;
        RECT  0.08 0.96 0.38 1.24 ;
        RECT  0.08 0.96 0.24 2.20 ;
        RECT  0.08 1.92 0.38 2.20 ;
        RECT  0.08 2.04 0.98 2.20 ;
        RECT  0.82 2.04 0.98 2.64 ;
        RECT  0.82 2.48 1.92 2.64 ;
        RECT  1.64 2.48 1.92 2.76 ;
        RECT  3.26 0.76 3.58 1.04 ;
        RECT  3.26 0.76 3.42 2.00 ;
        RECT  2.92 1.84 3.96 2.00 ;
        RECT  2.92 1.84 3.20 2.12 ;
        RECT  3.68 1.84 3.96 2.12 ;
        RECT  3.82 0.76 4.10 1.04 ;
        RECT  3.94 0.76 4.10 1.36 ;
        RECT  4.78 1.08 5.06 1.36 ;
        RECT  3.94 1.20 5.06 1.36 ;
        RECT  4.20 1.20 4.36 2.12 ;
        RECT  4.20 1.84 4.48 2.12 ;
        RECT  2.30 0.86 2.58 1.14 ;
        RECT  1.74 0.98 2.58 1.14 ;
        RECT  1.74 0.96 2.02 1.24 ;
        RECT  1.96 0.98 2.12 2.12 ;
        RECT  2.08 1.84 2.24 2.44 ;
        RECT  2.08 2.28 5.18 2.44 ;
        RECT  4.90 2.28 5.18 2.56 ;
        RECT  4.34 0.76 5.62 0.92 ;
        RECT  4.34 0.76 4.62 1.04 ;
        RECT  5.34 0.76 5.62 1.16 ;
        RECT  5.34 0.76 5.50 1.68 ;
        RECT  6.38 1.40 6.66 1.68 ;
        RECT  4.92 1.52 6.66 1.68 ;
        RECT  5.68 1.52 5.84 2.12 ;
        RECT  4.92 1.52 5.08 2.12 ;
        RECT  4.72 1.84 5.08 2.12 ;
        RECT  5.68 1.84 6.04 2.12 ;
        RECT  2.94 0.44 6.54 0.60 ;
        RECT  6.38 0.44 6.54 1.04 ;
        RECT  6.38 0.88 7.04 1.04 ;
        RECT  2.94 0.44 3.10 1.14 ;
        RECT  6.76 0.88 7.04 1.16 ;
        RECT  2.82 0.86 2.98 1.46 ;
        RECT  2.60 1.30 2.98 1.46 ;
        RECT  6.82 0.88 6.98 2.12 ;
        RECT  2.60 1.30 2.76 2.12 ;
        RECT  2.48 1.84 2.76 2.12 ;
        RECT  6.76 1.84 7.04 2.12 ;
        RECT  7.38 0.88 7.66 1.16 ;
        RECT  7.38 1.00 7.92 1.16 ;
        RECT  7.76 1.00 7.92 2.12 ;
        RECT  7.76 1.84 8.04 2.12 ;
        RECT  7.76 1.96 8.64 2.12 ;
        RECT  8.48 1.96 8.64 2.64 ;
        RECT  8.48 2.48 9.11 2.64 ;
        RECT  8.83 2.48 9.11 2.76 ;
        RECT  8.80 0.88 9.08 1.16 ;
        RECT  8.10 1.46 9.22 1.62 ;
        RECT  8.10 1.40 8.38 1.68 ;
        RECT  8.92 1.40 9.22 1.68 ;
        RECT  8.92 0.88 9.08 2.12 ;
        RECT  8.80 1.84 9.08 2.12 ;
    END
END DFFDSSP1V1_0

MACRO DFFDSP8V1_1
    CLASS CORE ;
    FOREIGN DFFDSP8V1_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 21.51  LAYER ME1  ;
        ANTENNADIFFAREA 11.20  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.56  LAYER ME1  ;
        ANTENNAMAXAREACAR 13.83  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.70 1.84 10.98 2.12 ;
        RECT  10.70 0.96 10.98 1.24 ;
        RECT  10.70 0.96 10.86 2.12 ;
        RECT  10.46 1.46 10.86 1.74 ;
        RECT  9.78 1.52 10.86 1.68 ;
        RECT  9.66 1.84 9.94 2.12 ;
        RECT  9.78 0.96 9.94 2.12 ;
        RECT  9.66 0.96 9.94 1.24 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 21.51  LAYER ME1  ;
        ANTENNADIFFAREA 11.40  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.56  LAYER ME1  ;
        ANTENNAMAXAREACAR 13.83  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.62 1.84 8.90 2.12 ;
        RECT  8.62 0.96 8.90 1.24 ;
        RECT  8.62 0.96 8.78 2.12 ;
        RECT  7.66 1.52 8.78 1.68 ;
        RECT  7.66 1.46 7.94 1.74 ;
        RECT  7.58 1.84 7.86 2.12 ;
        RECT  7.66 0.96 7.86 2.12 ;
        RECT  7.58 0.96 7.86 1.24 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.39 0.72 1.81 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.88 1.39 1.16 1.81 ;
        END
    END CK
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 11.60 0.28 ;
        RECT  11.22 0.64 11.50 0.92 ;
        RECT  11.28 -0.28 11.44 0.92 ;
        RECT  11.14 -0.28 11.44 0.32 ;
        RECT  10.18 0.64 10.46 0.92 ;
        RECT  10.24 -0.28 10.40 0.92 ;
        RECT  9.14 0.64 9.42 0.92 ;
        RECT  9.20 -0.28 9.36 0.92 ;
        RECT  8.10 0.64 8.38 0.92 ;
        RECT  8.16 -0.28 8.32 0.92 ;
        RECT  7.06 0.64 7.34 0.92 ;
        RECT  7.12 -0.28 7.28 0.92 ;
        RECT  6.06 0.96 6.34 1.24 ;
        RECT  6.16 -0.28 6.32 1.24 ;
        RECT  3.34 0.72 3.62 1.00 ;
        RECT  3.40 -0.28 3.56 1.00 ;
        RECT  0.62 0.68 0.90 0.96 ;
        RECT  0.68 -0.28 0.84 0.96 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 11.60 3.48 ;
        RECT  11.22 2.16 11.50 2.44 ;
        RECT  11.14 2.88 11.44 3.48 ;
        RECT  11.28 2.16 11.44 3.48 ;
        RECT  10.18 2.16 10.46 2.44 ;
        RECT  10.24 2.16 10.40 3.48 ;
        RECT  9.14 2.16 9.42 2.44 ;
        RECT  9.20 2.16 9.36 3.48 ;
        RECT  8.10 2.16 8.38 2.44 ;
        RECT  8.16 2.16 8.32 3.48 ;
        RECT  7.06 1.84 7.34 2.12 ;
        RECT  7.12 1.84 7.28 3.48 ;
        RECT  6.06 2.62 6.34 3.48 ;
        RECT  3.48 1.92 3.76 2.20 ;
        RECT  3.54 1.92 3.70 3.48 ;
        RECT  0.38 2.62 0.66 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  1.14 0.68 1.48 0.96 ;
        RECT  1.32 1.22 1.64 1.50 ;
        RECT  1.32 0.68 1.48 2.25 ;
        RECT  1.14 1.97 1.48 2.25 ;
        RECT  0.08 0.68 0.38 0.96 ;
        RECT  1.68 0.72 1.96 1.00 ;
        RECT  0.08 0.68 0.24 2.25 ;
        RECT  0.08 1.97 0.38 2.25 ;
        RECT  1.80 0.72 1.96 2.20 ;
        RECT  0.08 2.09 0.98 2.25 ;
        RECT  0.82 2.09 0.98 2.57 ;
        RECT  1.68 1.92 1.84 2.57 ;
        RECT  0.82 2.41 1.84 2.57 ;
        RECT  2.76 0.72 3.05 1.00 ;
        RECT  2.76 0.72 2.92 2.20 ;
        RECT  2.72 1.92 3.00 2.20 ;
        RECT  2.20 0.72 2.48 1.00 ;
        RECT  3.56 1.48 3.84 1.76 ;
        RECT  3.16 1.60 3.84 1.76 ;
        RECT  2.26 0.72 2.42 2.20 ;
        RECT  2.20 1.92 2.48 2.20 ;
        RECT  2.32 1.92 2.48 2.52 ;
        RECT  3.16 1.60 3.32 2.52 ;
        RECT  2.32 2.36 3.32 2.52 ;
        RECT  3.86 0.72 4.16 1.00 ;
        RECT  3.08 1.16 4.16 1.32 ;
        RECT  3.08 1.16 3.36 1.44 ;
        RECT  4.00 0.72 4.16 2.20 ;
        RECT  4.00 1.92 4.28 2.20 ;
        RECT  4.54 0.44 6.00 0.60 ;
        RECT  5.72 0.44 6.00 0.80 ;
        RECT  4.54 0.44 4.70 1.04 ;
        RECT  4.42 0.76 4.70 1.04 ;
        RECT  4.52 0.76 4.68 2.20 ;
        RECT  4.52 1.92 4.80 2.20 ;
        RECT  5.54 0.96 5.82 1.24 ;
        RECT  5.54 1.46 6.54 1.62 ;
        RECT  6.26 1.40 6.54 1.68 ;
        RECT  5.54 0.96 5.70 2.12 ;
        RECT  5.54 1.84 5.82 2.12 ;
        RECT  4.94 0.76 5.22 1.04 ;
        RECT  6.58 0.96 6.86 1.24 ;
        RECT  6.58 1.84 6.86 2.12 ;
        RECT  5.06 0.76 5.22 2.20 ;
        RECT  5.04 1.92 5.32 2.20 ;
        RECT  5.16 1.92 5.32 2.44 ;
        RECT  6.70 0.96 6.86 2.70 ;
        RECT  5.16 2.28 6.86 2.44 ;
        RECT  6.68 2.42 6.96 2.70 ;
    END
END DFFDSP8V1_1

MACRO DFFDSP8V1_0
    CLASS CORE ;
    FOREIGN DFFDSP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 22.67  LAYER ME1  ;
        ANTENNADIFFAREA 11.76  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.79  LAYER ME1  ;
        ANTENNAMAXAREACAR 12.66  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.36 1.84 11.64 2.12 ;
        RECT  11.36 0.96 11.64 1.24 ;
        RECT  11.36 0.96 11.52 2.12 ;
        RECT  10.06 1.46 11.52 1.62 ;
        RECT  10.32 1.84 10.60 2.12 ;
        RECT  10.32 0.96 10.60 1.24 ;
        RECT  10.32 0.96 10.48 2.12 ;
        RECT  10.06 1.46 10.48 1.74 ;
        END
    END Q
    PIN QB
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 22.67  LAYER ME1  ;
        ANTENNADIFFAREA 11.76  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.79  LAYER ME1  ;
        ANTENNAMAXAREACAR 12.66  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.28 1.84 9.56 2.12 ;
        RECT  9.28 0.96 9.56 1.24 ;
        RECT  9.34 0.96 9.50 2.12 ;
        RECT  8.36 1.46 9.50 1.62 ;
        RECT  8.36 1.46 8.74 1.74 ;
        RECT  8.24 1.84 8.52 2.12 ;
        RECT  8.36 0.96 8.52 2.12 ;
        RECT  8.24 0.96 8.52 1.24 ;
        END
    END QB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.46 1.39 0.74 1.81 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.66 1.34 1.94 1.76 ;
        END
    END D
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 12.40 0.28 ;
        RECT  11.94 -0.28 12.22 0.32 ;
        RECT  11.88 0.64 12.16 0.92 ;
        RECT  11.94 -0.28 12.10 0.92 ;
        RECT  10.84 0.64 11.12 0.92 ;
        RECT  10.90 -0.28 11.06 0.92 ;
        RECT  9.80 0.64 10.08 0.92 ;
        RECT  9.86 -0.28 10.02 0.92 ;
        RECT  8.76 0.64 9.04 0.92 ;
        RECT  8.82 -0.28 8.98 0.92 ;
        RECT  7.72 0.64 8.00 0.92 ;
        RECT  7.78 -0.28 7.94 0.92 ;
        RECT  6.72 0.96 7.00 1.24 ;
        RECT  6.82 -0.28 6.98 1.24 ;
        RECT  4.00 0.68 4.28 0.96 ;
        RECT  4.06 -0.28 4.22 0.96 ;
        RECT  1.64 0.68 1.92 0.96 ;
        RECT  1.70 -0.28 1.86 0.96 ;
        RECT  0.62 0.50 0.90 0.78 ;
        RECT  0.68 -0.28 0.84 0.78 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 12.40 3.48 ;
        RECT  11.94 2.88 12.22 3.48 ;
        RECT  11.88 2.16 12.16 2.44 ;
        RECT  11.94 2.16 12.10 3.48 ;
        RECT  10.84 2.16 11.12 2.44 ;
        RECT  10.90 2.16 11.06 3.48 ;
        RECT  9.80 2.16 10.08 2.44 ;
        RECT  9.86 2.16 10.02 3.48 ;
        RECT  8.76 2.16 9.04 2.44 ;
        RECT  8.82 2.16 8.98 3.48 ;
        RECT  7.72 1.84 8.00 2.12 ;
        RECT  7.78 1.84 7.94 3.48 ;
        RECT  6.72 2.62 7.00 3.48 ;
        RECT  4.00 1.92 4.28 2.20 ;
        RECT  4.06 1.92 4.22 3.48 ;
        RECT  1.76 1.92 1.92 3.48 ;
        RECT  1.64 1.92 1.92 2.20 ;
        RECT  0.62 1.97 0.90 2.25 ;
        RECT  0.68 1.97 0.84 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.08 0.50 0.38 0.78 ;
        RECT  0.08 1.00 1.16 1.16 ;
        RECT  0.88 0.94 1.16 1.22 ;
        RECT  0.08 0.50 0.24 2.25 ;
        RECT  0.08 1.97 0.38 2.25 ;
        RECT  1.14 0.50 1.48 0.78 ;
        RECT  1.14 1.97 1.48 2.25 ;
        RECT  1.32 0.50 1.48 2.70 ;
        RECT  1.32 2.42 1.60 2.70 ;
        RECT  2.16 0.68 2.44 0.96 ;
        RECT  2.22 0.68 2.38 2.20 ;
        RECT  2.16 1.92 2.44 2.20 ;
        RECT  2.68 0.68 2.96 0.96 ;
        RECT  2.74 0.68 2.90 2.20 ;
        RECT  2.68 1.92 2.96 2.20 ;
        RECT  2.80 1.92 2.96 2.70 ;
        RECT  3.34 2.42 3.62 2.70 ;
        RECT  2.80 2.54 3.62 2.70 ;
        RECT  3.34 0.68 3.62 0.96 ;
        RECT  3.40 0.68 3.56 2.20 ;
        RECT  3.34 1.92 3.62 2.20 ;
        RECT  4.52 0.68 4.80 0.96 ;
        RECT  3.86 1.44 4.74 1.60 ;
        RECT  3.86 1.38 4.14 1.66 ;
        RECT  4.58 0.68 4.74 2.20 ;
        RECT  4.52 1.92 4.80 2.20 ;
        RECT  5.20 0.44 6.66 0.60 ;
        RECT  6.38 0.44 6.66 0.80 ;
        RECT  5.20 0.44 5.36 1.04 ;
        RECT  5.08 0.76 5.36 1.04 ;
        RECT  5.10 0.76 5.26 2.20 ;
        RECT  5.04 1.92 5.32 2.20 ;
        RECT  6.20 0.96 6.48 1.24 ;
        RECT  6.20 1.46 7.19 1.62 ;
        RECT  6.91 1.40 7.19 1.68 ;
        RECT  6.20 0.96 6.36 2.12 ;
        RECT  6.20 1.84 6.48 2.12 ;
        RECT  5.60 0.76 5.88 1.04 ;
        RECT  7.24 0.96 7.52 1.24 ;
        RECT  7.36 0.96 7.52 2.12 ;
        RECT  5.62 0.76 5.78 2.20 ;
        RECT  5.56 1.92 5.84 2.20 ;
        RECT  5.68 1.92 5.84 2.44 ;
        RECT  7.24 1.84 7.40 2.44 ;
        RECT  5.68 2.28 7.62 2.44 ;
        RECT  7.34 2.28 7.62 2.71 ;
    END
END DFFDSP8V1_0

MACRO DFFDSP4V1_1
    CLASS CORE ;
    FOREIGN DFFDSP4V1_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 17.71  LAYER ME1  ;
        ANTENNADIFFAREA 8.66  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.98  LAYER ME1  ;
        ANTENNAMAXAREACAR 18.08  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.82 1.46 9.14 1.74 ;
        RECT  8.70 1.84 8.98 2.12 ;
        RECT  8.82 0.96 8.98 2.12 ;
        RECT  8.70 0.96 8.98 1.24 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 18.01  LAYER ME1  ;
        ANTENNADIFFAREA 8.66  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.98  LAYER ME1  ;
        ANTENNAMAXAREACAR 18.39  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.66 0.96 7.94 2.12 ;
        END
    END QB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.88 1.39 1.16 1.81 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.39 0.72 1.81 ;
        END
    END D
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 9.60 0.28 ;
        RECT  9.22 0.64 9.50 0.92 ;
        RECT  9.28 -0.28 9.44 0.92 ;
        RECT  9.14 -0.28 9.44 0.32 ;
        RECT  8.18 0.64 8.46 0.92 ;
        RECT  8.24 -0.28 8.40 0.92 ;
        RECT  7.14 0.64 7.42 0.92 ;
        RECT  7.20 -0.28 7.36 0.92 ;
        RECT  6.14 0.96 6.42 1.24 ;
        RECT  6.24 -0.28 6.40 1.24 ;
        RECT  3.36 0.72 3.64 1.00 ;
        RECT  3.42 -0.28 3.58 1.00 ;
        RECT  0.62 0.68 0.90 0.96 ;
        RECT  0.68 -0.28 0.84 0.96 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 9.60 3.48 ;
        RECT  9.22 2.16 9.50 2.44 ;
        RECT  9.14 2.88 9.44 3.48 ;
        RECT  9.28 2.16 9.44 3.48 ;
        RECT  8.18 2.16 8.46 2.44 ;
        RECT  8.24 2.16 8.40 3.48 ;
        RECT  7.14 1.84 7.42 2.12 ;
        RECT  7.20 1.84 7.36 3.48 ;
        RECT  6.14 2.62 6.42 3.48 ;
        RECT  3.48 1.92 3.76 2.20 ;
        RECT  3.54 1.92 3.70 3.48 ;
        RECT  0.38 2.62 0.66 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  1.14 0.68 1.48 0.96 ;
        RECT  1.32 1.22 1.64 1.50 ;
        RECT  1.32 0.68 1.48 2.25 ;
        RECT  1.14 1.97 1.48 2.25 ;
        RECT  0.08 0.68 0.38 0.96 ;
        RECT  1.68 0.72 1.96 1.00 ;
        RECT  0.08 0.68 0.24 2.25 ;
        RECT  0.08 1.97 0.38 2.25 ;
        RECT  1.80 0.72 1.96 2.20 ;
        RECT  0.08 2.09 0.98 2.25 ;
        RECT  0.82 2.09 0.98 2.57 ;
        RECT  1.68 1.92 1.84 2.57 ;
        RECT  0.82 2.41 1.84 2.57 ;
        RECT  2.76 0.72 3.07 1.00 ;
        RECT  2.76 0.72 2.92 2.20 ;
        RECT  2.72 1.92 3.00 2.20 ;
        RECT  2.20 0.72 2.48 1.00 ;
        RECT  3.56 1.48 3.84 1.76 ;
        RECT  3.16 1.60 3.84 1.76 ;
        RECT  2.26 0.72 2.42 2.20 ;
        RECT  2.20 1.92 2.48 2.20 ;
        RECT  2.32 1.92 2.48 2.52 ;
        RECT  3.16 1.60 3.32 2.52 ;
        RECT  2.32 2.36 3.32 2.52 ;
        RECT  3.88 0.72 4.16 1.00 ;
        RECT  3.08 1.16 4.16 1.32 ;
        RECT  3.08 1.16 3.36 1.44 ;
        RECT  4.00 0.72 4.16 2.20 ;
        RECT  4.00 1.92 4.28 2.20 ;
        RECT  4.62 0.44 6.08 0.60 ;
        RECT  5.80 0.44 6.08 0.80 ;
        RECT  4.62 0.44 4.78 1.04 ;
        RECT  4.50 0.76 4.78 1.04 ;
        RECT  4.58 0.76 4.74 2.20 ;
        RECT  4.52 1.92 4.80 2.20 ;
        RECT  5.62 0.96 5.90 1.24 ;
        RECT  5.62 1.46 6.62 1.62 ;
        RECT  6.34 1.40 6.62 1.68 ;
        RECT  5.62 0.96 5.78 2.12 ;
        RECT  5.62 1.84 5.90 2.12 ;
        RECT  5.02 0.76 5.30 1.04 ;
        RECT  6.66 0.96 6.94 1.24 ;
        RECT  6.66 1.84 6.94 2.12 ;
        RECT  5.10 0.76 5.26 2.20 ;
        RECT  5.04 1.92 5.32 2.20 ;
        RECT  5.16 1.92 5.32 2.44 ;
        RECT  6.78 0.96 6.94 2.70 ;
        RECT  5.16 2.28 6.94 2.44 ;
        RECT  6.76 2.42 7.04 2.70 ;
    END
END DFFDSP4V1_1

MACRO DFFDSP4V1_0
    CLASS CORE ;
    FOREIGN DFFDSP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 19.09  LAYER ME1  ;
        ANTENNADIFFAREA 9.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.21  LAYER ME1  ;
        ANTENNAMAXAREACAR 15.72  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.26 1.46 9.56 2.12 ;
        RECT  9.28 0.96 9.56 1.24 ;
        RECT  9.32 0.96 9.48 2.12 ;
        END
    END Q
    PIN QB
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 19.09  LAYER ME1  ;
        ANTENNADIFFAREA 9.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.21  LAYER ME1  ;
        ANTENNAMAXAREACAR 15.72  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.36 1.46 8.74 1.74 ;
        RECT  8.24 1.84 8.52 2.12 ;
        RECT  8.36 0.96 8.52 2.12 ;
        RECT  8.24 0.96 8.52 1.24 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.66 1.34 1.94 1.76 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.46 1.39 0.74 1.81 ;
        END
    END CK
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 10.40 3.48 ;
        RECT  9.86 2.88 10.22 3.48 ;
        RECT  9.80 2.16 10.08 2.44 ;
        RECT  9.86 2.16 10.02 3.48 ;
        RECT  8.76 2.16 9.04 2.44 ;
        RECT  8.82 2.16 8.98 3.48 ;
        RECT  7.72 1.87 8.00 2.15 ;
        RECT  7.78 1.87 7.94 3.48 ;
        RECT  6.72 2.62 7.00 3.48 ;
        RECT  4.00 1.92 4.28 2.20 ;
        RECT  4.06 1.92 4.22 3.48 ;
        RECT  1.76 1.92 1.92 3.48 ;
        RECT  1.64 1.92 1.92 2.20 ;
        RECT  0.62 1.97 0.90 2.25 ;
        RECT  0.68 1.97 0.84 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 10.40 0.28 ;
        RECT  9.86 -0.28 10.22 0.32 ;
        RECT  9.80 0.64 10.08 0.92 ;
        RECT  9.86 -0.28 10.02 0.92 ;
        RECT  8.76 0.64 9.04 0.92 ;
        RECT  8.82 -0.28 8.98 0.92 ;
        RECT  7.72 0.64 8.00 0.92 ;
        RECT  7.78 -0.28 7.94 0.92 ;
        RECT  6.72 0.96 7.00 1.24 ;
        RECT  6.82 -0.28 6.98 1.24 ;
        RECT  4.00 0.68 4.28 0.96 ;
        RECT  4.06 -0.28 4.22 0.96 ;
        RECT  1.64 0.68 1.92 0.96 ;
        RECT  1.70 -0.28 1.86 0.96 ;
        RECT  0.62 0.50 0.90 0.78 ;
        RECT  0.68 -0.28 0.84 0.78 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.08 0.50 0.38 0.78 ;
        RECT  0.08 1.00 1.16 1.16 ;
        RECT  0.88 0.94 1.16 1.22 ;
        RECT  0.08 0.50 0.24 2.25 ;
        RECT  0.08 1.97 0.38 2.25 ;
        RECT  1.14 0.50 1.48 0.78 ;
        RECT  1.14 1.97 1.48 2.25 ;
        RECT  1.32 0.50 1.48 2.70 ;
        RECT  1.32 2.42 1.60 2.70 ;
        RECT  2.16 0.68 2.44 0.96 ;
        RECT  2.22 0.68 2.38 2.20 ;
        RECT  2.16 1.92 2.44 2.20 ;
        RECT  2.68 0.68 2.96 0.96 ;
        RECT  2.74 0.68 2.90 2.20 ;
        RECT  2.68 1.92 2.96 2.20 ;
        RECT  2.80 1.92 2.96 2.70 ;
        RECT  3.34 2.42 3.62 2.70 ;
        RECT  2.80 2.54 3.62 2.70 ;
        RECT  3.34 0.68 3.62 0.96 ;
        RECT  3.40 0.68 3.56 2.20 ;
        RECT  3.34 1.92 3.62 2.20 ;
        RECT  4.52 0.68 4.80 0.96 ;
        RECT  3.86 1.44 4.74 1.60 ;
        RECT  3.86 1.38 4.14 1.66 ;
        RECT  4.58 0.68 4.74 2.20 ;
        RECT  4.52 1.92 4.80 2.20 ;
        RECT  5.20 0.44 6.66 0.60 ;
        RECT  6.38 0.44 6.66 0.80 ;
        RECT  5.20 0.44 5.36 1.04 ;
        RECT  5.08 0.76 5.36 1.04 ;
        RECT  5.10 0.76 5.26 2.20 ;
        RECT  5.04 1.92 5.32 2.20 ;
        RECT  6.20 0.96 6.48 1.24 ;
        RECT  6.20 1.46 7.19 1.62 ;
        RECT  6.91 1.40 7.19 1.68 ;
        RECT  6.20 0.96 6.36 2.12 ;
        RECT  6.20 1.84 6.48 2.12 ;
        RECT  5.60 0.76 5.88 1.04 ;
        RECT  7.24 0.96 7.52 1.24 ;
        RECT  7.36 0.96 7.52 2.12 ;
        RECT  5.62 0.76 5.78 2.20 ;
        RECT  5.56 1.92 5.84 2.20 ;
        RECT  5.68 1.92 5.84 2.44 ;
        RECT  7.24 1.84 7.40 2.44 ;
        RECT  5.68 2.28 7.62 2.44 ;
        RECT  7.34 2.28 7.62 2.71 ;
    END
END DFFDSP4V1_0

MACRO DFFDSP2V1_1
    CLASS CORE ;
    FOREIGN DFFDSP2V1_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.39 0.72 1.81 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.88 1.39 1.16 1.81 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 16.19  LAYER ME1  ;
        ANTENNADIFFAREA 7.45  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.69  LAYER ME1  ;
        ANTENNAMAXAREACAR 23.42  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.26 1.46 7.54 1.74 ;
        RECT  7.16 1.84 7.44 2.12 ;
        RECT  7.26 0.96 7.44 2.12 ;
        RECT  7.16 0.96 7.44 1.24 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 16.48  LAYER ME1  ;
        ANTENNADIFFAREA 7.45  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.69  LAYER ME1  ;
        ANTENNAMAXAREACAR 23.84  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.32 1.46 8.72 1.74 ;
        RECT  8.20 1.84 8.48 2.12 ;
        RECT  8.32 0.96 8.48 2.12 ;
        RECT  8.20 0.96 8.48 1.24 ;
        END
    END Q
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 8.80 3.48 ;
        RECT  8.34 2.88 8.62 3.48 ;
        RECT  7.68 2.16 7.96 2.44 ;
        RECT  7.74 2.16 7.90 3.48 ;
        RECT  6.16 2.62 6.44 3.48 ;
        RECT  3.48 1.92 3.76 2.20 ;
        RECT  3.54 1.92 3.70 3.48 ;
        RECT  0.38 2.62 0.66 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 8.80 0.28 ;
        RECT  8.34 -0.28 8.62 0.32 ;
        RECT  7.68 0.64 7.96 0.92 ;
        RECT  7.74 -0.28 7.90 0.92 ;
        RECT  6.16 0.96 6.44 1.24 ;
        RECT  6.26 -0.28 6.42 1.24 ;
        RECT  3.36 0.72 3.64 1.00 ;
        RECT  3.42 -0.28 3.58 1.00 ;
        RECT  0.62 0.68 0.90 0.96 ;
        RECT  0.68 -0.28 0.84 0.96 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  1.14 0.68 1.48 0.96 ;
        RECT  1.32 1.22 1.64 1.50 ;
        RECT  1.32 0.68 1.48 2.25 ;
        RECT  1.14 1.97 1.48 2.25 ;
        RECT  0.08 0.68 0.38 0.96 ;
        RECT  1.68 0.72 1.96 1.00 ;
        RECT  0.08 0.68 0.24 2.25 ;
        RECT  0.08 1.97 0.38 2.25 ;
        RECT  1.80 0.72 1.96 2.20 ;
        RECT  0.08 2.09 0.98 2.25 ;
        RECT  0.82 2.09 0.98 2.57 ;
        RECT  1.68 1.92 1.84 2.57 ;
        RECT  0.82 2.41 1.84 2.57 ;
        RECT  2.76 0.72 3.07 1.00 ;
        RECT  2.76 0.72 2.92 2.20 ;
        RECT  2.72 1.92 3.00 2.20 ;
        RECT  2.20 0.72 2.48 1.00 ;
        RECT  3.56 1.48 3.84 1.76 ;
        RECT  3.16 1.60 3.84 1.76 ;
        RECT  2.26 0.72 2.42 2.20 ;
        RECT  2.20 1.92 2.48 2.20 ;
        RECT  2.32 1.92 2.48 2.52 ;
        RECT  3.16 1.60 3.32 2.52 ;
        RECT  2.32 2.36 3.32 2.52 ;
        RECT  3.88 0.72 4.16 1.00 ;
        RECT  3.08 1.16 4.16 1.32 ;
        RECT  3.08 1.16 3.36 1.44 ;
        RECT  4.00 0.72 4.16 2.20 ;
        RECT  4.00 1.92 4.28 2.20 ;
        RECT  4.64 0.44 6.10 0.60 ;
        RECT  5.82 0.44 6.10 0.80 ;
        RECT  4.64 0.44 4.80 1.04 ;
        RECT  4.52 0.76 4.80 1.04 ;
        RECT  4.58 0.76 4.74 2.20 ;
        RECT  4.52 1.92 4.80 2.20 ;
        RECT  5.64 0.96 5.92 1.24 ;
        RECT  5.64 1.46 6.64 1.62 ;
        RECT  6.36 1.40 6.64 1.68 ;
        RECT  5.64 0.96 5.80 2.12 ;
        RECT  5.64 1.84 5.92 2.12 ;
        RECT  5.04 0.76 5.32 1.04 ;
        RECT  6.68 0.96 6.96 1.24 ;
        RECT  6.68 1.84 6.96 2.12 ;
        RECT  5.10 0.76 5.26 2.20 ;
        RECT  5.04 1.92 5.32 2.20 ;
        RECT  5.16 1.92 5.32 2.44 ;
        RECT  6.80 0.96 6.96 2.70 ;
        RECT  5.16 2.28 6.96 2.44 ;
        RECT  6.78 2.42 7.06 2.70 ;
    END
END DFFDSP2V1_1

MACRO DFFDSP2V1_0
    CLASS CORE ;
    FOREIGN DFFDSP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 17.03  LAYER ME1  ;
        ANTENNADIFFAREA 7.65  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.93  LAYER ME1  ;
        ANTENNAMAXAREACAR 18.38  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.76 1.84 9.08 2.12 ;
        RECT  8.92 0.96 9.08 2.12 ;
        RECT  8.76 0.96 9.08 1.24 ;
        END
    END Q
    PIN QB
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 16.78  LAYER ME1  ;
        ANTENNADIFFAREA 7.65  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.93  LAYER ME1  ;
        ANTENNAMAXAREACAR 18.11  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.72 1.84 8.00 2.12 ;
        RECT  7.72 0.96 8.00 1.24 ;
        RECT  7.72 0.96 7.88 2.12 ;
        END
    END QB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.46 1.39 0.74 1.81 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.66 1.34 1.94 1.76 ;
        END
    END D
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 9.20 0.28 ;
        RECT  8.74 -0.28 9.02 0.32 ;
        RECT  8.24 0.64 8.52 0.92 ;
        RECT  8.30 -0.28 8.46 0.92 ;
        RECT  6.72 0.96 7.00 1.24 ;
        RECT  6.82 -0.28 6.98 1.24 ;
        RECT  4.00 0.68 4.28 0.96 ;
        RECT  4.06 -0.28 4.22 0.96 ;
        RECT  1.64 0.68 1.92 0.96 ;
        RECT  1.70 -0.28 1.86 0.96 ;
        RECT  0.62 0.50 0.90 0.78 ;
        RECT  0.68 -0.28 0.84 0.78 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 9.20 3.48 ;
        RECT  8.74 2.88 9.02 3.48 ;
        RECT  8.24 2.16 8.52 2.44 ;
        RECT  8.30 2.16 8.46 3.48 ;
        RECT  6.72 2.62 7.00 3.48 ;
        RECT  4.00 1.92 4.28 2.20 ;
        RECT  4.06 1.92 4.22 3.48 ;
        RECT  1.76 1.92 1.92 3.48 ;
        RECT  1.64 1.92 1.92 2.20 ;
        RECT  0.62 1.97 0.90 2.25 ;
        RECT  0.68 1.97 0.84 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.08 0.50 0.38 0.78 ;
        RECT  0.08 1.00 1.16 1.16 ;
        RECT  0.88 0.94 1.16 1.22 ;
        RECT  0.08 0.50 0.24 2.25 ;
        RECT  0.08 1.97 0.38 2.25 ;
        RECT  1.14 0.50 1.48 0.78 ;
        RECT  1.14 1.97 1.48 2.25 ;
        RECT  1.32 0.50 1.48 2.70 ;
        RECT  1.32 2.42 1.60 2.70 ;
        RECT  2.16 0.68 2.44 0.96 ;
        RECT  2.22 0.68 2.38 2.20 ;
        RECT  2.16 1.92 2.44 2.20 ;
        RECT  2.68 0.68 2.96 0.96 ;
        RECT  2.74 0.68 2.90 2.20 ;
        RECT  2.68 1.92 2.96 2.20 ;
        RECT  2.80 1.92 2.96 2.70 ;
        RECT  3.34 2.42 3.62 2.70 ;
        RECT  2.80 2.54 3.62 2.70 ;
        RECT  3.34 0.68 3.62 0.96 ;
        RECT  3.40 0.68 3.56 2.20 ;
        RECT  3.34 1.92 3.62 2.20 ;
        RECT  4.52 0.68 4.80 0.96 ;
        RECT  3.86 1.44 4.74 1.60 ;
        RECT  3.86 1.38 4.14 1.66 ;
        RECT  4.58 0.68 4.74 2.20 ;
        RECT  4.52 1.92 4.80 2.20 ;
        RECT  5.20 0.44 6.66 0.60 ;
        RECT  6.38 0.44 6.66 0.80 ;
        RECT  5.20 0.44 5.36 1.04 ;
        RECT  5.08 0.76 5.36 1.04 ;
        RECT  5.10 0.76 5.26 2.20 ;
        RECT  5.04 1.92 5.32 2.20 ;
        RECT  6.20 0.96 6.48 1.24 ;
        RECT  6.20 1.46 7.19 1.62 ;
        RECT  6.91 1.40 7.19 1.68 ;
        RECT  6.20 0.96 6.36 2.12 ;
        RECT  6.20 1.84 6.48 2.12 ;
        RECT  5.60 0.76 5.88 1.04 ;
        RECT  7.24 0.96 7.52 1.24 ;
        RECT  7.36 0.96 7.52 2.12 ;
        RECT  5.62 0.76 5.78 2.20 ;
        RECT  5.56 1.92 5.84 2.20 ;
        RECT  5.68 1.92 5.84 2.44 ;
        RECT  7.24 1.84 7.40 2.44 ;
        RECT  5.68 2.28 7.62 2.44 ;
        RECT  7.34 2.28 7.62 2.71 ;
    END
END DFFDSP2V1_0

MACRO DFFDSP1V1_1
    CLASS CORE ;
    FOREIGN DFFDSP1V1_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 16.58  LAYER ME1  ;
        ANTENNADIFFAREA 6.76  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.54  LAYER ME1  ;
        ANTENNAMAXAREACAR 30.84  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.32 1.46 8.72 1.74 ;
        RECT  8.20 1.84 8.48 2.12 ;
        RECT  8.32 0.96 8.48 2.12 ;
        RECT  8.20 0.96 8.48 1.24 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 16.29  LAYER ME1  ;
        ANTENNADIFFAREA 6.76  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.54  LAYER ME1  ;
        ANTENNAMAXAREACAR 30.30  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.26 1.46 7.54 1.74 ;
        RECT  7.16 1.84 7.44 2.12 ;
        RECT  7.26 0.96 7.44 2.12 ;
        RECT  7.16 0.96 7.44 1.24 ;
        END
    END QB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.88 1.39 1.16 1.81 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.39 0.72 1.81 ;
        END
    END D
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 8.80 0.28 ;
        RECT  8.34 -0.28 8.62 0.32 ;
        RECT  7.68 0.96 7.96 1.24 ;
        RECT  7.74 -0.28 7.90 1.24 ;
        RECT  6.16 0.96 6.44 1.24 ;
        RECT  6.26 -0.28 6.42 1.24 ;
        RECT  3.36 0.72 3.64 1.00 ;
        RECT  3.42 -0.28 3.58 1.00 ;
        RECT  0.62 0.68 0.90 0.96 ;
        RECT  0.68 -0.28 0.84 0.96 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 8.80 3.48 ;
        RECT  8.34 2.88 8.62 3.48 ;
        RECT  7.68 1.84 7.96 2.12 ;
        RECT  7.74 1.84 7.90 3.48 ;
        RECT  6.16 2.62 6.44 3.48 ;
        RECT  3.48 1.92 3.76 2.20 ;
        RECT  3.54 1.92 3.70 3.48 ;
        RECT  0.38 2.62 0.66 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  1.14 0.68 1.48 0.96 ;
        RECT  1.32 1.22 1.64 1.50 ;
        RECT  1.32 0.68 1.48 2.25 ;
        RECT  1.14 1.97 1.48 2.25 ;
        RECT  0.08 0.68 0.38 0.96 ;
        RECT  1.68 0.72 1.96 1.00 ;
        RECT  0.08 0.68 0.24 2.25 ;
        RECT  0.08 1.97 0.38 2.25 ;
        RECT  1.80 0.72 1.96 2.20 ;
        RECT  0.08 2.09 0.98 2.25 ;
        RECT  0.82 2.09 0.98 2.57 ;
        RECT  1.68 1.92 1.84 2.57 ;
        RECT  0.82 2.41 1.84 2.57 ;
        RECT  2.76 0.72 3.07 1.00 ;
        RECT  2.76 0.72 2.92 2.20 ;
        RECT  2.72 1.92 3.00 2.20 ;
        RECT  2.20 0.72 2.48 1.00 ;
        RECT  3.56 1.48 3.84 1.76 ;
        RECT  3.16 1.60 3.84 1.76 ;
        RECT  2.26 0.72 2.42 2.20 ;
        RECT  2.20 1.92 2.48 2.20 ;
        RECT  2.32 1.92 2.48 2.52 ;
        RECT  3.16 1.60 3.32 2.52 ;
        RECT  2.32 2.36 3.32 2.52 ;
        RECT  3.88 0.72 4.16 1.00 ;
        RECT  3.08 1.16 4.16 1.32 ;
        RECT  3.08 1.16 3.36 1.44 ;
        RECT  4.00 0.72 4.16 2.20 ;
        RECT  4.00 1.92 4.28 2.20 ;
        RECT  4.64 0.44 6.10 0.60 ;
        RECT  5.82 0.44 6.10 0.80 ;
        RECT  4.64 0.44 4.80 1.04 ;
        RECT  4.52 0.76 4.80 1.04 ;
        RECT  4.58 0.76 4.74 2.20 ;
        RECT  4.52 1.92 4.80 2.20 ;
        RECT  5.64 0.96 5.92 1.24 ;
        RECT  5.64 1.46 6.64 1.62 ;
        RECT  6.36 1.40 6.64 1.68 ;
        RECT  5.64 0.96 5.80 2.12 ;
        RECT  5.64 1.84 5.92 2.12 ;
        RECT  5.04 0.76 5.32 1.04 ;
        RECT  6.68 0.96 6.96 1.24 ;
        RECT  6.68 1.84 6.96 2.12 ;
        RECT  5.10 0.76 5.26 2.20 ;
        RECT  5.04 1.92 5.32 2.20 ;
        RECT  5.16 1.92 5.32 2.44 ;
        RECT  6.80 0.96 6.96 2.44 ;
        RECT  5.16 2.28 7.10 2.44 ;
        RECT  6.82 2.28 7.10 2.62 ;
    END
END DFFDSP1V1_1

MACRO DFFDSP1V1_0
    CLASS CORE ;
    FOREIGN DFFDSP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.66 1.34 1.94 1.76 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.46 1.39 0.74 1.81 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 17.14  LAYER ME1  ;
        ANTENNADIFFAREA 6.96  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.77  LAYER ME1  ;
        ANTENNAMAXAREACAR 22.18  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.76 1.84 9.08 2.12 ;
        RECT  8.92 0.96 9.08 2.12 ;
        RECT  8.76 0.96 9.08 1.24 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 16.89  LAYER ME1  ;
        ANTENNADIFFAREA 6.96  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.77  LAYER ME1  ;
        ANTENNAMAXAREACAR 21.85  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.72 1.84 8.00 2.12 ;
        RECT  7.72 0.96 8.00 1.24 ;
        RECT  7.72 0.96 7.88 2.12 ;
        END
    END QB
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 9.20 3.48 ;
        RECT  8.74 2.88 9.02 3.48 ;
        RECT  8.24 1.84 8.52 2.12 ;
        RECT  8.30 1.84 8.46 3.48 ;
        RECT  6.72 2.62 7.00 3.48 ;
        RECT  4.00 1.92 4.28 2.20 ;
        RECT  4.06 1.92 4.22 3.48 ;
        RECT  1.64 1.92 1.92 2.20 ;
        RECT  1.72 1.92 1.88 3.48 ;
        RECT  0.62 1.97 0.90 2.25 ;
        RECT  0.68 1.97 0.84 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 9.20 0.28 ;
        RECT  8.74 -0.28 9.02 0.32 ;
        RECT  8.24 0.96 8.52 1.24 ;
        RECT  8.30 -0.28 8.46 1.24 ;
        RECT  6.72 0.96 7.00 1.24 ;
        RECT  6.82 -0.28 6.98 1.24 ;
        RECT  4.00 0.68 4.28 0.96 ;
        RECT  4.06 -0.28 4.22 0.96 ;
        RECT  1.64 0.68 1.92 0.96 ;
        RECT  1.70 -0.28 1.86 0.96 ;
        RECT  0.62 0.50 0.90 0.78 ;
        RECT  0.68 -0.28 0.84 0.78 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.08 0.50 0.38 0.78 ;
        RECT  0.08 1.00 1.16 1.16 ;
        RECT  0.88 0.94 1.16 1.22 ;
        RECT  0.08 0.50 0.24 2.25 ;
        RECT  0.08 1.97 0.38 2.25 ;
        RECT  1.14 0.50 1.48 0.78 ;
        RECT  1.14 1.97 1.48 2.25 ;
        RECT  1.32 0.50 1.48 2.70 ;
        RECT  1.28 2.42 1.56 2.70 ;
        RECT  2.16 0.68 2.44 0.96 ;
        RECT  2.22 0.68 2.38 2.20 ;
        RECT  2.16 1.92 2.44 2.20 ;
        RECT  2.68 0.68 2.96 0.96 ;
        RECT  2.68 1.92 2.96 2.20 ;
        RECT  2.74 0.68 2.90 2.70 ;
        RECT  3.34 2.42 3.62 2.70 ;
        RECT  2.74 2.54 3.62 2.70 ;
        RECT  3.34 0.68 3.62 0.96 ;
        RECT  3.40 0.68 3.56 2.20 ;
        RECT  3.34 1.92 3.62 2.20 ;
        RECT  4.52 0.68 4.80 0.96 ;
        RECT  3.86 1.44 4.74 1.60 ;
        RECT  3.86 1.38 4.14 1.66 ;
        RECT  4.58 0.68 4.74 2.20 ;
        RECT  4.52 1.92 4.80 2.20 ;
        RECT  5.20 0.44 6.66 0.60 ;
        RECT  6.38 0.44 6.66 0.80 ;
        RECT  5.20 0.44 5.36 1.04 ;
        RECT  5.08 0.76 5.36 1.04 ;
        RECT  5.10 0.76 5.26 2.20 ;
        RECT  5.04 1.92 5.32 2.20 ;
        RECT  6.20 0.96 6.48 1.24 ;
        RECT  6.20 1.46 7.20 1.62 ;
        RECT  6.92 1.40 7.20 1.68 ;
        RECT  6.20 0.96 6.36 2.12 ;
        RECT  6.20 1.84 6.48 2.12 ;
        RECT  5.60 0.76 5.88 1.04 ;
        RECT  7.24 0.96 7.52 1.24 ;
        RECT  7.24 1.84 7.52 2.12 ;
        RECT  5.62 0.76 5.78 2.20 ;
        RECT  5.56 1.92 5.84 2.20 ;
        RECT  5.68 1.92 5.84 2.44 ;
        RECT  7.36 0.96 7.52 2.44 ;
        RECT  5.68 2.28 7.76 2.44 ;
        RECT  7.48 2.28 7.76 2.62 ;
    END
END DFFDSP1V1_0

MACRO DFFDRZSP8V1_0
    CLASS CORE ;
    FOREIGN DFFDRZSP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 30.30  LAYER ME1  ;
        ANTENNADIFFAREA 14.81  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.62  LAYER ME1  ;
        ANTENNAMAXAREACAR 18.68  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.91 1.90 15.19 2.50 ;
        RECT  14.91 0.64 15.19 1.24 ;
        RECT  14.91 0.64 15.07 2.50 ;
        RECT  13.99 1.52 15.07 1.68 ;
        RECT  13.99 1.46 14.34 1.74 ;
        RECT  13.87 1.90 14.15 2.50 ;
        RECT  13.99 0.64 14.15 2.50 ;
        RECT  13.87 0.64 14.15 1.24 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 30.30  LAYER ME1  ;
        ANTENNADIFFAREA 14.56  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.62  LAYER ME1  ;
        ANTENNAMAXAREACAR 18.68  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.83 1.90 13.11 2.50 ;
        RECT  12.83 0.64 13.11 1.24 ;
        RECT  12.83 0.64 12.99 2.50 ;
        RECT  11.66 1.52 12.99 1.68 ;
        RECT  11.79 1.90 12.07 2.50 ;
        RECT  11.79 0.64 12.07 1.24 ;
        RECT  11.79 0.64 11.95 2.50 ;
        RECT  11.66 1.46 11.95 1.74 ;
        END
    END Q
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.22 1.40 9.60 1.68 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.21 1.40 3.53 1.76 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.87  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 12.90  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.06 1.46 2.34 1.74 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.81 2.23 2.25 ;
        RECT  1.95 0.81 2.23 1.09 ;
        END
    END TD
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END SEL
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.20  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.83  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.81 1.19 2.25 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  0.91 0.81 1.19 1.09 ;
        END
    END D
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 16.00 0.28 ;
        RECT  15.49 -0.28 15.82 0.32 ;
        RECT  15.43 0.64 15.71 1.24 ;
        RECT  15.49 -0.28 15.65 1.24 ;
        RECT  14.39 0.64 14.67 1.24 ;
        RECT  14.45 -0.28 14.61 1.24 ;
        RECT  13.35 0.64 13.63 1.24 ;
        RECT  13.41 -0.28 13.57 1.24 ;
        RECT  12.31 0.64 12.59 1.24 ;
        RECT  12.37 -0.28 12.53 1.24 ;
        RECT  11.27 0.64 11.55 1.24 ;
        RECT  11.33 -0.28 11.49 1.24 ;
        RECT  10.27 0.88 10.55 1.16 ;
        RECT  10.33 -0.28 10.49 1.16 ;
        RECT  7.29 -0.28 7.57 0.72 ;
        RECT  2.71 -0.28 2.99 0.68 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 16.00 3.48 ;
        RECT  15.49 2.88 15.82 3.48 ;
        RECT  15.43 1.90 15.71 2.50 ;
        RECT  15.49 1.90 15.65 3.48 ;
        RECT  14.39 1.90 14.67 2.50 ;
        RECT  14.45 1.90 14.61 3.48 ;
        RECT  13.35 1.90 13.63 2.50 ;
        RECT  13.41 1.90 13.57 3.48 ;
        RECT  12.31 1.90 12.59 2.50 ;
        RECT  12.37 1.90 12.53 3.48 ;
        RECT  11.27 1.90 11.55 2.50 ;
        RECT  11.33 1.90 11.49 3.48 ;
        RECT  10.27 1.84 10.55 2.12 ;
        RECT  10.33 1.84 10.49 3.48 ;
        RECT  9.23 1.84 9.51 2.12 ;
        RECT  9.29 1.84 9.45 3.48 ;
        RECT  8.39 1.84 8.55 3.48 ;
        RECT  8.19 1.84 8.55 2.12 ;
        RECT  2.71 2.52 2.99 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  1.55 1.97 1.71 2.57 ;
        RECT  1.55 2.41 2.37 2.57 ;
        RECT  2.09 2.41 2.37 2.69 ;
        RECT  3.47 0.96 3.85 1.24 ;
        RECT  3.69 1.46 3.97 1.74 ;
        RECT  3.69 0.96 3.85 2.20 ;
        RECT  3.47 1.92 3.85 2.20 ;
        RECT  4.07 0.44 4.35 0.72 ;
        RECT  3.15 0.56 4.35 0.72 ;
        RECT  3.15 0.56 3.31 1.12 ;
        RECT  2.43 0.96 3.31 1.12 ;
        RECT  2.43 0.96 2.71 1.24 ;
        RECT  2.50 0.96 2.66 2.20 ;
        RECT  2.43 1.92 2.71 2.20 ;
        RECT  2.43 2.04 3.31 2.20 ;
        RECT  3.15 2.04 3.31 2.64 ;
        RECT  3.15 2.48 4.35 2.64 ;
        RECT  4.07 2.48 4.35 2.76 ;
        RECT  5.67 0.88 5.95 1.16 ;
        RECT  5.67 0.88 5.83 2.12 ;
        RECT  5.45 1.84 5.83 2.12 ;
        RECT  6.15 1.84 6.43 2.12 ;
        RECT  5.45 1.96 6.43 2.12 ;
        RECT  6.85 0.44 7.13 0.72 ;
        RECT  6.31 0.56 7.13 0.72 ;
        RECT  6.19 0.88 6.47 1.16 ;
        RECT  6.31 0.56 6.47 1.68 ;
        RECT  6.31 1.52 6.75 1.68 ;
        RECT  6.59 1.52 6.75 2.12 ;
        RECT  6.59 1.84 6.95 2.12 ;
        RECT  4.63 0.87 4.91 1.15 ;
        RECT  4.07 0.99 4.91 1.15 ;
        RECT  4.07 0.96 4.35 1.24 ;
        RECT  4.19 0.96 4.35 2.12 ;
        RECT  4.19 1.84 4.47 2.12 ;
        RECT  4.19 1.96 4.77 2.12 ;
        RECT  4.61 1.96 4.77 2.76 ;
        RECT  7.95 2.42 8.23 2.76 ;
        RECT  4.61 2.60 8.23 2.76 ;
        RECT  8.15 0.50 8.43 0.78 ;
        RECT  6.71 0.88 6.99 1.20 ;
        RECT  7.33 0.92 7.61 1.20 ;
        RECT  8.15 0.50 8.31 1.20 ;
        RECT  6.71 1.04 8.31 1.20 ;
        RECT  7.11 1.04 7.27 2.12 ;
        RECT  7.11 1.84 7.47 2.12 ;
        RECT  5.13 0.87 5.43 1.15 ;
        RECT  8.81 0.92 9.09 1.20 ;
        RECT  7.63 1.52 8.97 1.68 ;
        RECT  8.81 0.92 8.97 2.12 ;
        RECT  5.01 1.84 5.29 2.12 ;
        RECT  8.71 1.84 8.99 2.12 ;
        RECT  5.13 0.87 5.29 2.44 ;
        RECT  7.63 1.52 7.79 2.44 ;
        RECT  5.13 2.28 7.79 2.44 ;
        RECT  9.37 0.88 9.65 1.16 ;
        RECT  9.37 1.00 9.92 1.16 ;
        RECT  9.76 1.46 10.75 1.62 ;
        RECT  10.47 1.40 10.75 1.68 ;
        RECT  9.76 1.00 9.92 2.12 ;
        RECT  9.75 1.84 10.03 2.12 ;
        RECT  10.79 0.88 11.07 1.16 ;
        RECT  10.79 1.84 11.07 2.12 ;
        RECT  10.91 0.88 11.07 2.76 ;
        RECT  10.82 2.48 11.10 2.76 ;
    END
END DFFDRZSP8V1_0

MACRO DFFDRZSP4V1_0
    CLASS CORE ;
    FOREIGN DFFDRZSP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.20  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.83  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.81 1.19 2.25 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  0.91 0.81 1.19 1.09 ;
        END
    END D
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END SEL
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.87  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 12.90  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.06 1.46 2.34 1.74 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.81 2.23 2.25 ;
        RECT  1.95 0.81 2.23 1.09 ;
        END
    END TD
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.21 1.40 3.53 1.76 ;
        END
    END CK
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.22 1.40 9.60 1.68 ;
        END
    END RB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 26.05  LAYER ME1  ;
        ANTENNADIFFAREA 11.52  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.05  LAYER ME1  ;
        ANTENNAMAXAREACAR 24.89  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.79 1.90 12.07 2.50 ;
        RECT  11.79 0.64 12.07 1.24 ;
        RECT  11.79 0.64 11.95 2.50 ;
        RECT  11.66 1.46 11.95 1.74 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 26.05  LAYER ME1  ;
        ANTENNADIFFAREA 11.77  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.05  LAYER ME1  ;
        ANTENNAMAXAREACAR 24.89  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.86 1.46 13.14 1.74 ;
        RECT  12.83 1.90 13.11 2.50 ;
        RECT  12.86 0.64 13.11 2.50 ;
        RECT  12.83 0.64 13.11 1.24 ;
        END
    END QB
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 14.00 3.48 ;
        RECT  13.41 2.88 13.82 3.48 ;
        RECT  13.35 1.90 13.63 2.50 ;
        RECT  13.41 1.90 13.57 3.48 ;
        RECT  12.31 1.90 12.59 2.50 ;
        RECT  12.37 1.90 12.53 3.48 ;
        RECT  11.27 1.90 11.55 2.50 ;
        RECT  11.33 1.90 11.49 3.48 ;
        RECT  10.27 1.84 10.55 2.12 ;
        RECT  10.33 1.84 10.49 3.48 ;
        RECT  9.23 1.84 9.51 2.12 ;
        RECT  9.29 1.84 9.45 3.48 ;
        RECT  8.39 1.84 8.55 3.48 ;
        RECT  8.19 1.84 8.55 2.12 ;
        RECT  2.71 2.52 2.99 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 14.00 0.28 ;
        RECT  13.41 -0.28 13.82 0.32 ;
        RECT  13.35 0.64 13.63 1.24 ;
        RECT  13.41 -0.28 13.57 1.24 ;
        RECT  12.31 0.64 12.59 1.24 ;
        RECT  12.37 -0.28 12.53 1.24 ;
        RECT  11.27 0.64 11.55 1.24 ;
        RECT  11.33 -0.28 11.49 1.24 ;
        RECT  10.27 0.88 10.55 1.16 ;
        RECT  10.33 -0.28 10.49 1.16 ;
        RECT  7.29 -0.28 7.57 0.72 ;
        RECT  2.71 -0.28 2.99 0.68 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  1.55 1.97 1.71 2.57 ;
        RECT  1.55 2.41 2.37 2.57 ;
        RECT  2.09 2.41 2.37 2.69 ;
        RECT  3.47 0.96 3.85 1.24 ;
        RECT  3.69 1.46 3.97 1.74 ;
        RECT  3.69 0.96 3.85 2.20 ;
        RECT  3.47 1.92 3.85 2.20 ;
        RECT  4.07 0.44 4.35 0.72 ;
        RECT  3.15 0.56 4.35 0.72 ;
        RECT  3.15 0.56 3.31 1.12 ;
        RECT  2.43 0.96 3.31 1.12 ;
        RECT  2.43 0.96 2.71 1.24 ;
        RECT  2.50 0.96 2.66 2.20 ;
        RECT  2.43 1.92 2.71 2.20 ;
        RECT  2.43 2.04 3.31 2.20 ;
        RECT  3.15 2.04 3.31 2.64 ;
        RECT  3.15 2.48 4.35 2.64 ;
        RECT  4.07 2.48 4.35 2.76 ;
        RECT  5.67 0.88 5.95 1.16 ;
        RECT  5.67 0.88 5.83 2.12 ;
        RECT  5.45 1.84 5.83 2.12 ;
        RECT  6.15 1.84 6.43 2.12 ;
        RECT  5.45 1.96 6.43 2.12 ;
        RECT  6.85 0.44 7.13 0.72 ;
        RECT  6.31 0.56 7.13 0.72 ;
        RECT  6.19 0.88 6.47 1.16 ;
        RECT  6.31 0.56 6.47 1.68 ;
        RECT  6.31 1.52 6.75 1.68 ;
        RECT  6.59 1.52 6.75 2.12 ;
        RECT  6.59 1.84 6.95 2.12 ;
        RECT  4.63 0.87 4.91 1.15 ;
        RECT  4.07 0.99 4.91 1.15 ;
        RECT  4.07 0.96 4.35 1.24 ;
        RECT  4.19 0.96 4.35 2.12 ;
        RECT  4.19 1.84 4.47 2.12 ;
        RECT  4.19 1.96 4.77 2.12 ;
        RECT  4.61 1.96 4.77 2.76 ;
        RECT  7.95 2.42 8.23 2.76 ;
        RECT  4.61 2.60 8.23 2.76 ;
        RECT  8.15 0.50 8.43 0.78 ;
        RECT  6.71 0.88 6.99 1.20 ;
        RECT  7.33 0.92 7.61 1.20 ;
        RECT  8.15 0.50 8.31 1.20 ;
        RECT  6.71 1.04 8.31 1.20 ;
        RECT  7.11 1.04 7.27 2.12 ;
        RECT  7.11 1.84 7.47 2.12 ;
        RECT  5.13 0.87 5.43 1.15 ;
        RECT  8.81 0.92 9.09 1.20 ;
        RECT  7.63 1.52 8.97 1.68 ;
        RECT  8.81 0.92 8.97 2.12 ;
        RECT  5.01 1.84 5.29 2.12 ;
        RECT  8.71 1.84 8.99 2.12 ;
        RECT  5.13 0.87 5.29 2.44 ;
        RECT  7.63 1.52 7.79 2.44 ;
        RECT  5.13 2.28 7.79 2.44 ;
        RECT  9.37 0.88 9.65 1.16 ;
        RECT  9.37 1.00 9.92 1.16 ;
        RECT  9.76 1.46 10.75 1.62 ;
        RECT  10.47 1.40 10.75 1.68 ;
        RECT  9.76 1.00 9.92 2.12 ;
        RECT  9.75 1.84 10.03 2.12 ;
        RECT  10.79 0.88 11.07 1.16 ;
        RECT  10.79 1.84 11.07 2.12 ;
        RECT  10.91 0.88 11.07 2.76 ;
        RECT  10.82 2.48 11.10 2.76 ;
    END
END DFFDRZSP4V1_0

MACRO DFFDRZSP2V1_0
    CLASS CORE ;
    FOREIGN DFFDRZSP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 23.79  LAYER ME1  ;
        ANTENNADIFFAREA 10.19  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.76  LAYER ME1  ;
        ANTENNAMAXAREACAR 31.37  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.43 1.46 12.72 1.74 ;
        RECT  12.31 1.90 12.59 2.50 ;
        RECT  12.43 0.64 12.59 2.50 ;
        RECT  12.31 0.64 12.59 1.24 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 23.79  LAYER ME1  ;
        ANTENNADIFFAREA 10.19  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.76  LAYER ME1  ;
        ANTENNAMAXAREACAR 31.37  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.27 1.90 11.55 2.50 ;
        RECT  11.27 0.64 11.55 1.24 ;
        RECT  11.27 0.64 11.54 2.50 ;
        RECT  11.26 1.46 11.54 1.74 ;
        END
    END Q
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.22 1.40 9.60 1.68 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.21 1.40 3.53 1.76 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.87  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 12.90  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.06 1.46 2.34 1.74 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.81 2.23 2.25 ;
        RECT  1.95 0.81 2.23 1.09 ;
        END
    END TD
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END SEL
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.20  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.83  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.81 1.19 2.25 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  0.91 0.81 1.19 1.09 ;
        END
    END D
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 12.80 0.28 ;
        RECT  12.34 -0.28 12.62 0.32 ;
        RECT  11.79 0.64 12.07 1.24 ;
        RECT  11.85 -0.28 12.01 1.24 ;
        RECT  10.27 0.88 10.55 1.16 ;
        RECT  10.33 -0.28 10.49 1.16 ;
        RECT  7.29 -0.28 7.57 0.72 ;
        RECT  2.71 -0.28 2.99 0.68 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 12.80 3.48 ;
        RECT  12.34 2.88 12.62 3.48 ;
        RECT  11.79 1.90 12.07 2.50 ;
        RECT  11.85 1.90 12.01 3.48 ;
        RECT  10.27 1.84 10.55 2.12 ;
        RECT  10.33 1.84 10.49 3.48 ;
        RECT  9.23 1.84 9.51 2.12 ;
        RECT  9.29 1.84 9.45 3.48 ;
        RECT  8.39 1.84 8.55 3.48 ;
        RECT  8.19 1.84 8.55 2.12 ;
        RECT  2.71 2.52 2.99 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  1.55 1.97 1.71 2.57 ;
        RECT  1.55 2.41 2.37 2.57 ;
        RECT  2.09 2.41 2.37 2.69 ;
        RECT  3.47 0.96 3.85 1.24 ;
        RECT  3.69 1.46 3.97 1.74 ;
        RECT  3.69 0.96 3.85 2.20 ;
        RECT  3.47 1.92 3.85 2.20 ;
        RECT  4.07 0.44 4.35 0.72 ;
        RECT  3.15 0.56 4.35 0.72 ;
        RECT  3.15 0.56 3.31 1.12 ;
        RECT  2.43 0.96 3.31 1.12 ;
        RECT  2.43 0.96 2.71 1.24 ;
        RECT  2.50 0.96 2.66 2.20 ;
        RECT  2.43 1.92 2.71 2.20 ;
        RECT  2.43 2.04 3.31 2.20 ;
        RECT  3.15 2.04 3.31 2.64 ;
        RECT  3.15 2.48 4.35 2.64 ;
        RECT  4.07 2.48 4.35 2.76 ;
        RECT  5.67 0.88 5.95 1.16 ;
        RECT  5.67 0.88 5.83 2.12 ;
        RECT  5.45 1.84 5.83 2.12 ;
        RECT  6.15 1.84 6.43 2.12 ;
        RECT  5.45 1.96 6.43 2.12 ;
        RECT  6.85 0.44 7.13 0.72 ;
        RECT  6.31 0.56 7.13 0.72 ;
        RECT  6.19 0.88 6.47 1.16 ;
        RECT  6.31 0.56 6.47 1.68 ;
        RECT  6.31 1.52 6.75 1.68 ;
        RECT  6.59 1.52 6.75 2.12 ;
        RECT  6.59 1.84 6.95 2.12 ;
        RECT  4.63 0.87 4.91 1.15 ;
        RECT  4.07 0.99 4.91 1.15 ;
        RECT  4.07 0.96 4.35 1.24 ;
        RECT  4.19 0.96 4.35 2.12 ;
        RECT  4.19 1.84 4.47 2.12 ;
        RECT  4.19 1.96 4.77 2.12 ;
        RECT  4.61 1.96 4.77 2.76 ;
        RECT  7.95 2.42 8.23 2.76 ;
        RECT  4.61 2.60 8.23 2.76 ;
        RECT  8.15 0.50 8.43 0.78 ;
        RECT  6.71 0.88 6.99 1.20 ;
        RECT  7.33 0.92 7.61 1.20 ;
        RECT  8.15 0.50 8.31 1.20 ;
        RECT  6.71 1.04 8.31 1.20 ;
        RECT  7.11 1.04 7.27 2.12 ;
        RECT  7.11 1.84 7.47 2.12 ;
        RECT  5.13 0.87 5.43 1.15 ;
        RECT  8.81 0.92 9.09 1.20 ;
        RECT  7.63 1.52 8.97 1.68 ;
        RECT  8.81 0.92 8.97 2.12 ;
        RECT  5.01 1.84 5.29 2.12 ;
        RECT  8.71 1.84 8.99 2.12 ;
        RECT  5.13 0.87 5.29 2.44 ;
        RECT  7.63 1.52 7.79 2.44 ;
        RECT  5.13 2.28 7.79 2.44 ;
        RECT  9.37 0.88 9.65 1.16 ;
        RECT  9.37 1.00 9.92 1.16 ;
        RECT  9.76 1.46 10.75 1.62 ;
        RECT  10.47 1.40 10.75 1.68 ;
        RECT  9.76 1.00 9.92 2.12 ;
        RECT  9.75 1.84 10.03 2.12 ;
        RECT  10.79 0.88 11.07 1.16 ;
        RECT  10.79 1.84 11.07 2.12 ;
        RECT  10.91 0.88 11.07 2.76 ;
        RECT  10.82 2.48 11.10 2.76 ;
    END
END DFFDRZSP2V1_0

MACRO DFFDRZSP1V1_0
    CLASS CORE ;
    FOREIGN DFFDRZSP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 23.06  LAYER ME1  ;
        ANTENNADIFFAREA 9.50  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.60  LAYER ME1  ;
        ANTENNAMAXAREACAR 38.14  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.43 1.46 12.72 1.74 ;
        RECT  12.31 1.90 12.59 2.18 ;
        RECT  12.43 0.88 12.59 2.18 ;
        RECT  12.31 0.88 12.59 1.16 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 23.38  LAYER ME1  ;
        ANTENNADIFFAREA 9.50  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.60  LAYER ME1  ;
        ANTENNAMAXAREACAR 38.65  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.27 1.90 11.55 2.18 ;
        RECT  11.27 0.88 11.55 1.16 ;
        RECT  11.27 0.88 11.54 2.18 ;
        RECT  11.26 1.46 11.54 1.74 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.20  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.83  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.81 1.19 2.25 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  0.91 0.81 1.19 1.09 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.21 1.40 3.53 1.76 ;
        END
    END CK
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.22 1.40 9.60 1.68 ;
        END
    END RB
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.87  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 12.90  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.06 1.46 2.34 1.74 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.81 2.23 2.25 ;
        RECT  1.95 0.81 2.23 1.09 ;
        END
    END TD
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END SEL
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 12.80 0.28 ;
        RECT  12.34 -0.28 12.62 0.32 ;
        RECT  11.79 0.88 12.07 1.16 ;
        RECT  11.85 -0.28 12.01 1.16 ;
        RECT  10.27 0.88 10.55 1.16 ;
        RECT  10.33 -0.28 10.49 1.16 ;
        RECT  7.29 -0.28 7.57 0.72 ;
        RECT  2.71 -0.28 2.99 0.68 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 12.80 3.48 ;
        RECT  12.34 2.88 12.62 3.48 ;
        RECT  11.79 1.90 12.07 2.18 ;
        RECT  11.85 1.90 12.01 3.48 ;
        RECT  10.27 1.84 10.55 2.12 ;
        RECT  10.33 1.84 10.49 3.48 ;
        RECT  9.23 1.84 9.51 2.12 ;
        RECT  9.29 1.84 9.45 3.48 ;
        RECT  8.39 1.84 8.55 3.48 ;
        RECT  8.19 1.84 8.55 2.12 ;
        RECT  2.71 2.52 2.99 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  1.55 1.97 1.71 2.57 ;
        RECT  1.55 2.41 2.37 2.57 ;
        RECT  2.09 2.41 2.37 2.69 ;
        RECT  3.47 0.96 3.85 1.24 ;
        RECT  3.69 1.46 3.97 1.74 ;
        RECT  3.69 0.96 3.85 2.20 ;
        RECT  3.47 1.92 3.85 2.20 ;
        RECT  4.07 0.44 4.35 0.72 ;
        RECT  3.15 0.56 4.35 0.72 ;
        RECT  3.15 0.56 3.31 1.12 ;
        RECT  2.43 0.96 3.31 1.12 ;
        RECT  2.43 0.96 2.71 1.24 ;
        RECT  2.50 0.96 2.66 2.20 ;
        RECT  2.43 1.92 2.71 2.20 ;
        RECT  2.43 2.04 3.31 2.20 ;
        RECT  3.15 2.04 3.31 2.64 ;
        RECT  3.15 2.48 4.35 2.64 ;
        RECT  4.07 2.48 4.35 2.76 ;
        RECT  5.67 0.88 5.95 1.16 ;
        RECT  5.67 0.88 5.83 2.12 ;
        RECT  5.45 1.84 5.83 2.12 ;
        RECT  6.15 1.84 6.43 2.12 ;
        RECT  5.45 1.96 6.43 2.12 ;
        RECT  6.85 0.44 7.13 0.72 ;
        RECT  6.31 0.56 7.13 0.72 ;
        RECT  6.19 0.88 6.47 1.16 ;
        RECT  6.31 0.56 6.47 1.68 ;
        RECT  6.31 1.52 6.75 1.68 ;
        RECT  6.59 1.52 6.75 2.12 ;
        RECT  6.59 1.84 6.95 2.12 ;
        RECT  4.63 0.87 4.91 1.15 ;
        RECT  4.07 0.99 4.91 1.15 ;
        RECT  4.07 0.96 4.35 1.24 ;
        RECT  4.19 0.96 4.35 2.12 ;
        RECT  4.19 1.84 4.47 2.12 ;
        RECT  4.19 1.96 4.77 2.12 ;
        RECT  4.61 1.96 4.77 2.76 ;
        RECT  7.95 2.42 8.23 2.76 ;
        RECT  4.61 2.60 8.23 2.76 ;
        RECT  8.15 0.50 8.43 0.78 ;
        RECT  6.71 0.88 6.99 1.20 ;
        RECT  7.33 0.92 7.61 1.20 ;
        RECT  8.15 0.50 8.31 1.20 ;
        RECT  6.71 1.04 8.31 1.20 ;
        RECT  7.11 1.04 7.27 2.12 ;
        RECT  7.11 1.84 7.47 2.12 ;
        RECT  5.13 0.87 5.43 1.15 ;
        RECT  8.81 0.92 9.09 1.20 ;
        RECT  7.63 1.52 8.97 1.68 ;
        RECT  8.81 0.92 8.97 2.12 ;
        RECT  5.01 1.84 5.29 2.12 ;
        RECT  8.71 1.84 8.99 2.12 ;
        RECT  5.13 0.87 5.29 2.44 ;
        RECT  7.63 1.52 7.79 2.44 ;
        RECT  5.13 2.28 7.79 2.44 ;
        RECT  9.37 0.88 9.65 1.16 ;
        RECT  9.37 1.00 9.92 1.16 ;
        RECT  9.76 1.46 10.75 1.62 ;
        RECT  10.47 1.40 10.75 1.68 ;
        RECT  9.76 1.00 9.92 2.12 ;
        RECT  9.75 1.84 10.03 2.12 ;
        RECT  10.79 0.88 11.07 1.16 ;
        RECT  10.79 1.84 11.07 2.12 ;
        RECT  10.91 0.88 11.07 2.76 ;
        RECT  10.82 2.48 11.10 2.76 ;
    END
END DFFDRZSP1V1_0

MACRO DFFDRSZSP8V1_0
    CLASS CORE ;
    FOREIGN DFFDRSZSP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 17.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 32.94  LAYER ME1  ;
        ANTENNADIFFAREA 15.94  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.62  LAYER ME1  ;
        ANTENNAMAXAREACAR 20.30  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.47 1.90 14.75 2.50 ;
        RECT  14.47 0.64 14.75 1.24 ;
        RECT  14.47 0.64 14.63 2.50 ;
        RECT  13.55 1.52 14.63 1.68 ;
        RECT  13.55 1.46 13.94 1.74 ;
        RECT  13.43 1.90 13.71 2.50 ;
        RECT  13.55 0.64 13.71 2.50 ;
        RECT  13.43 0.64 13.71 1.24 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.66 0.44 11.94 0.94 ;
        RECT  11.45 0.44 11.94 0.72 ;
        END
    END SB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.99 1.40 10.41 1.68 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.24 1.40 3.54 1.76 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.20  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.83  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.81 1.19 2.25 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  0.91 0.81 1.19 1.09 ;
        END
    END D
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END SEL
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.87  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 12.90  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.06 1.46 2.34 1.74 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.81 2.23 2.25 ;
        RECT  1.95 0.81 2.23 1.09 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 32.94  LAYER ME1  ;
        ANTENNADIFFAREA 16.18  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.62  LAYER ME1  ;
        ANTENNAMAXAREACAR 20.30  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  16.55 1.90 16.83 2.50 ;
        RECT  16.55 0.64 16.83 1.24 ;
        RECT  16.55 0.64 16.71 2.50 ;
        RECT  15.63 1.52 16.71 1.68 ;
        RECT  15.63 1.46 15.95 1.74 ;
        RECT  15.51 1.90 15.79 2.50 ;
        RECT  15.63 0.64 15.79 2.50 ;
        RECT  15.51 0.64 15.79 1.24 ;
        END
    END QB
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 17.60 0.28 ;
        RECT  17.13 -0.28 17.42 0.32 ;
        RECT  17.07 0.64 17.35 1.24 ;
        RECT  17.13 -0.28 17.29 1.24 ;
        RECT  16.03 0.64 16.31 1.24 ;
        RECT  16.09 -0.28 16.25 1.24 ;
        RECT  14.99 0.64 15.27 1.24 ;
        RECT  15.05 -0.28 15.21 1.24 ;
        RECT  13.95 0.64 14.23 1.24 ;
        RECT  14.01 -0.28 14.17 1.24 ;
        RECT  12.91 0.64 13.19 1.24 ;
        RECT  12.97 -0.28 13.13 1.24 ;
        RECT  11.08 0.88 11.43 1.16 ;
        RECT  11.08 -0.28 11.24 1.16 ;
        RECT  8.69 -0.28 8.97 0.68 ;
        RECT  2.71 -0.28 2.99 0.68 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 17.60 3.48 ;
        RECT  17.13 2.88 17.42 3.48 ;
        RECT  17.07 1.90 17.35 2.50 ;
        RECT  17.13 1.90 17.29 3.48 ;
        RECT  16.03 1.90 16.31 2.50 ;
        RECT  16.09 1.90 16.25 3.48 ;
        RECT  14.99 1.90 15.27 2.50 ;
        RECT  15.05 1.90 15.21 3.48 ;
        RECT  13.95 1.90 14.23 2.50 ;
        RECT  14.01 1.90 14.17 3.48 ;
        RECT  12.91 1.90 13.19 2.50 ;
        RECT  12.97 1.90 13.13 3.48 ;
        RECT  12.31 2.40 12.59 3.48 ;
        RECT  11.09 1.84 11.37 2.12 ;
        RECT  11.15 1.84 11.31 3.48 ;
        RECT  10.05 1.84 10.33 2.12 ;
        RECT  10.11 1.84 10.27 3.48 ;
        RECT  8.77 1.96 9.29 2.12 ;
        RECT  9.01 1.84 9.29 2.12 ;
        RECT  8.65 2.52 8.93 3.48 ;
        RECT  8.77 1.96 8.93 3.48 ;
        RECT  2.71 2.52 2.99 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  1.55 1.97 1.71 2.57 ;
        RECT  1.55 2.41 2.37 2.57 ;
        RECT  2.09 2.41 2.37 2.69 ;
        RECT  3.47 0.96 3.86 1.24 ;
        RECT  3.70 1.46 4.02 1.74 ;
        RECT  3.70 0.96 3.86 2.20 ;
        RECT  3.47 1.92 3.86 2.20 ;
        RECT  4.07 0.44 4.35 0.72 ;
        RECT  3.15 0.56 4.35 0.72 ;
        RECT  3.15 0.56 3.31 1.12 ;
        RECT  2.43 0.96 3.31 1.12 ;
        RECT  2.43 0.96 2.71 1.24 ;
        RECT  2.50 0.96 2.66 2.20 ;
        RECT  2.43 1.92 2.71 2.20 ;
        RECT  2.43 2.04 3.31 2.20 ;
        RECT  3.15 2.04 3.31 2.64 ;
        RECT  3.15 2.48 4.25 2.64 ;
        RECT  3.97 2.48 4.25 2.76 ;
        RECT  5.59 0.88 5.91 1.16 ;
        RECT  5.59 0.88 5.75 2.00 ;
        RECT  5.25 1.84 6.23 2.00 ;
        RECT  5.25 1.84 5.53 2.12 ;
        RECT  5.95 1.84 6.23 2.12 ;
        RECT  6.15 0.88 6.43 1.16 ;
        RECT  6.27 0.88 6.43 1.58 ;
        RECT  7.11 1.14 7.39 1.58 ;
        RECT  6.27 1.42 7.39 1.58 ;
        RECT  6.39 1.42 6.55 2.12 ;
        RECT  6.39 1.84 6.75 2.12 ;
        RECT  4.75 0.50 8.15 0.66 ;
        RECT  7.87 0.50 8.15 0.78 ;
        RECT  4.63 0.86 4.91 1.14 ;
        RECT  4.75 0.50 4.91 1.14 ;
        RECT  4.07 0.98 4.91 1.14 ;
        RECT  4.07 0.96 4.35 1.24 ;
        RECT  4.29 0.98 4.45 2.12 ;
        RECT  4.29 1.84 4.57 2.12 ;
        RECT  9.13 0.50 9.41 0.78 ;
        RECT  6.67 0.82 7.71 0.98 ;
        RECT  6.67 0.82 6.95 1.16 ;
        RECT  9.13 0.50 9.29 1.16 ;
        RECT  7.55 1.00 9.29 1.16 ;
        RECT  7.55 0.96 7.91 1.24 ;
        RECT  7.85 1.00 8.01 2.12 ;
        RECT  6.99 1.84 7.27 2.12 ;
        RECT  7.85 1.84 8.19 2.12 ;
        RECT  6.99 1.96 8.19 2.12 ;
        RECT  5.07 0.86 5.43 1.14 ;
        RECT  9.67 0.96 10.11 1.24 ;
        RECT  5.07 0.86 5.23 1.48 ;
        RECT  8.35 1.52 9.83 1.68 ;
        RECT  4.81 1.84 5.09 2.12 ;
        RECT  9.67 0.96 9.83 2.12 ;
        RECT  9.53 1.84 9.83 2.12 ;
        RECT  4.93 1.32 5.09 2.44 ;
        RECT  8.35 1.52 8.51 2.44 ;
        RECT  4.93 2.28 8.51 2.44 ;
        RECT  10.31 0.88 10.73 1.16 ;
        RECT  10.57 1.46 12.11 1.62 ;
        RECT  11.83 1.40 12.11 1.68 ;
        RECT  10.57 0.88 10.73 2.12 ;
        RECT  10.57 1.84 10.85 2.12 ;
        RECT  12.11 0.88 12.47 1.16 ;
        RECT  12.31 0.88 12.47 2.16 ;
        RECT  12.31 1.88 12.59 2.16 ;
        RECT  11.82 2.00 12.59 2.16 ;
        RECT  11.82 2.00 11.98 2.76 ;
        RECT  11.70 2.48 11.98 2.76 ;
    END
END DFFDRSZSP8V1_0

MACRO DFFDRSZSP4V1_0
    CLASS CORE ;
    FOREIGN DFFDRSZSP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 28.75  LAYER ME1  ;
        ANTENNADIFFAREA 13.14  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.05  LAYER ME1  ;
        ANTENNAMAXAREACAR 27.48  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.47 1.90 14.75 2.50 ;
        RECT  14.47 0.64 14.75 1.24 ;
        RECT  14.47 0.64 14.74 2.50 ;
        RECT  14.46 1.46 14.74 1.74 ;
        END
    END QB
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.87  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 12.90  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.06 1.46 2.34 1.74 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.81 2.23 2.25 ;
        RECT  1.95 0.81 2.23 1.09 ;
        END
    END TD
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END SEL
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.20  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.83  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.81 1.19 2.25 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  0.91 0.81 1.19 1.09 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.24 1.40 3.54 1.76 ;
        END
    END CK
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.99 1.40 10.41 1.68 ;
        END
    END RB
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.66 0.44 11.94 0.94 ;
        RECT  11.45 0.44 11.94 0.72 ;
        END
    END SB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 28.75  LAYER ME1  ;
        ANTENNADIFFAREA 12.90  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.05  LAYER ME1  ;
        ANTENNAMAXAREACAR 27.48  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.55 1.46 13.94 1.74 ;
        RECT  13.43 1.90 13.71 2.50 ;
        RECT  13.55 0.64 13.71 2.50 ;
        RECT  13.43 0.64 13.71 1.24 ;
        END
    END Q
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 15.60 3.48 ;
        RECT  15.05 2.88 15.42 3.48 ;
        RECT  14.99 1.90 15.27 2.50 ;
        RECT  15.05 1.90 15.21 3.48 ;
        RECT  13.95 1.90 14.23 2.50 ;
        RECT  14.01 1.90 14.17 3.48 ;
        RECT  12.91 1.90 13.19 2.50 ;
        RECT  12.97 1.90 13.13 3.48 ;
        RECT  12.31 2.40 12.59 3.48 ;
        RECT  11.09 1.84 11.37 2.12 ;
        RECT  11.15 1.84 11.31 3.48 ;
        RECT  10.05 1.84 10.33 2.12 ;
        RECT  10.11 1.84 10.27 3.48 ;
        RECT  8.77 1.96 9.29 2.12 ;
        RECT  9.01 1.84 9.29 2.12 ;
        RECT  8.65 2.52 8.93 3.48 ;
        RECT  8.77 1.96 8.93 3.48 ;
        RECT  2.71 2.52 2.99 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 15.60 0.28 ;
        RECT  15.05 -0.28 15.42 0.32 ;
        RECT  14.99 0.64 15.27 1.24 ;
        RECT  15.05 -0.28 15.21 1.24 ;
        RECT  13.95 0.64 14.23 1.24 ;
        RECT  14.01 -0.28 14.17 1.24 ;
        RECT  12.91 0.64 13.19 1.24 ;
        RECT  12.97 -0.28 13.13 1.24 ;
        RECT  11.08 0.88 11.43 1.16 ;
        RECT  11.08 -0.28 11.24 1.16 ;
        RECT  8.69 -0.28 8.97 0.68 ;
        RECT  2.71 -0.28 2.99 0.68 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  1.55 1.97 1.71 2.57 ;
        RECT  1.55 2.41 2.37 2.57 ;
        RECT  2.09 2.41 2.37 2.69 ;
        RECT  3.47 0.96 3.86 1.24 ;
        RECT  3.70 1.46 4.02 1.74 ;
        RECT  3.70 0.96 3.86 2.20 ;
        RECT  3.47 1.92 3.86 2.20 ;
        RECT  4.07 0.44 4.35 0.72 ;
        RECT  3.15 0.56 4.35 0.72 ;
        RECT  3.15 0.56 3.31 1.12 ;
        RECT  2.43 0.96 3.31 1.12 ;
        RECT  2.43 0.96 2.71 1.24 ;
        RECT  2.50 0.96 2.66 2.20 ;
        RECT  2.43 1.92 2.71 2.20 ;
        RECT  2.43 2.04 3.31 2.20 ;
        RECT  3.15 2.04 3.31 2.64 ;
        RECT  3.15 2.48 4.25 2.64 ;
        RECT  3.97 2.48 4.25 2.76 ;
        RECT  5.59 0.88 5.91 1.16 ;
        RECT  5.59 0.88 5.75 2.00 ;
        RECT  5.25 1.84 6.23 2.00 ;
        RECT  5.25 1.84 5.53 2.12 ;
        RECT  5.95 1.84 6.23 2.12 ;
        RECT  6.15 0.88 6.43 1.16 ;
        RECT  6.27 0.88 6.43 1.58 ;
        RECT  7.11 1.14 7.39 1.58 ;
        RECT  6.27 1.42 7.39 1.58 ;
        RECT  6.39 1.42 6.55 2.12 ;
        RECT  6.39 1.84 6.75 2.12 ;
        RECT  4.75 0.50 8.15 0.66 ;
        RECT  7.87 0.50 8.15 0.78 ;
        RECT  4.63 0.86 4.91 1.14 ;
        RECT  4.75 0.50 4.91 1.14 ;
        RECT  4.07 0.98 4.91 1.14 ;
        RECT  4.07 0.96 4.35 1.24 ;
        RECT  4.29 0.98 4.45 2.12 ;
        RECT  4.29 1.84 4.57 2.12 ;
        RECT  9.13 0.50 9.41 0.78 ;
        RECT  6.67 0.82 7.71 0.98 ;
        RECT  6.67 0.82 6.95 1.16 ;
        RECT  9.13 0.50 9.29 1.16 ;
        RECT  7.55 1.00 9.29 1.16 ;
        RECT  7.55 0.96 7.91 1.24 ;
        RECT  7.85 1.00 8.01 2.12 ;
        RECT  6.99 1.84 7.27 2.12 ;
        RECT  7.85 1.84 8.19 2.12 ;
        RECT  6.99 1.96 8.19 2.12 ;
        RECT  5.07 0.86 5.43 1.14 ;
        RECT  9.67 0.96 10.11 1.24 ;
        RECT  5.07 0.86 5.23 1.48 ;
        RECT  8.35 1.52 9.83 1.68 ;
        RECT  4.81 1.84 5.09 2.12 ;
        RECT  9.67 0.96 9.83 2.12 ;
        RECT  9.53 1.84 9.83 2.12 ;
        RECT  4.93 1.32 5.09 2.44 ;
        RECT  8.35 1.52 8.51 2.44 ;
        RECT  4.93 2.28 8.51 2.44 ;
        RECT  10.31 0.88 10.73 1.16 ;
        RECT  10.57 1.46 12.11 1.62 ;
        RECT  11.83 1.40 12.11 1.68 ;
        RECT  10.57 0.88 10.73 2.12 ;
        RECT  10.57 1.84 10.85 2.12 ;
        RECT  12.11 0.88 12.47 1.16 ;
        RECT  12.31 0.88 12.47 2.16 ;
        RECT  12.31 1.88 12.59 2.16 ;
        RECT  11.82 2.00 12.59 2.16 ;
        RECT  11.82 2.00 11.98 2.76 ;
        RECT  11.70 2.48 11.98 2.76 ;
    END
END DFFDRSZSP4V1_0

MACRO DFFDRSZSP2V1_0
    CLASS CORE ;
    FOREIGN DFFDRSZSP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 26.44  LAYER ME1  ;
        ANTENNADIFFAREA 11.56  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.76  LAYER ME1  ;
        ANTENNAMAXAREACAR 34.87  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.06 1.46 14.32 1.74 ;
        RECT  13.95 1.89 14.23 2.49 ;
        RECT  14.06 0.64 14.23 2.49 ;
        RECT  13.95 0.64 14.23 1.24 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 26.44  LAYER ME1  ;
        ANTENNADIFFAREA 11.56  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.76  LAYER ME1  ;
        ANTENNAMAXAREACAR 34.87  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.91 1.89 13.19 2.49 ;
        RECT  12.91 0.64 13.19 1.24 ;
        RECT  12.91 0.64 13.14 2.49 ;
        RECT  12.85 1.46 13.14 1.74 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.66 0.44 11.94 0.94 ;
        RECT  11.45 0.44 11.94 0.72 ;
        END
    END SB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.99 1.40 10.41 1.68 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.24 1.40 3.54 1.76 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.20  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.83  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.81 1.19 2.25 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  0.91 0.81 1.19 1.09 ;
        END
    END D
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END SEL
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.87  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 12.90  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.06 1.46 2.34 1.74 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.81 2.23 2.25 ;
        RECT  1.95 0.81 2.23 1.09 ;
        END
    END TD
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 14.40 0.28 ;
        RECT  13.94 -0.28 14.22 0.32 ;
        RECT  13.43 0.64 13.71 1.24 ;
        RECT  13.49 -0.28 13.65 1.24 ;
        RECT  11.08 0.88 11.43 1.16 ;
        RECT  11.08 -0.28 11.24 1.16 ;
        RECT  8.69 -0.28 8.97 0.68 ;
        RECT  2.71 -0.28 2.99 0.68 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 14.40 3.48 ;
        RECT  13.94 2.88 14.22 3.48 ;
        RECT  13.43 1.89 13.71 2.49 ;
        RECT  13.49 1.89 13.65 3.48 ;
        RECT  12.31 2.40 12.59 3.48 ;
        RECT  11.09 1.84 11.37 2.12 ;
        RECT  11.15 1.84 11.31 3.48 ;
        RECT  10.05 1.84 10.33 2.12 ;
        RECT  10.11 1.84 10.27 3.48 ;
        RECT  8.77 1.96 9.29 2.12 ;
        RECT  9.01 1.84 9.29 2.12 ;
        RECT  8.65 2.52 8.93 3.48 ;
        RECT  8.77 1.96 8.93 3.48 ;
        RECT  2.71 2.52 2.99 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  1.55 1.97 1.71 2.57 ;
        RECT  1.55 2.41 2.37 2.57 ;
        RECT  2.09 2.41 2.37 2.69 ;
        RECT  3.47 0.96 3.86 1.24 ;
        RECT  3.70 1.46 4.02 1.74 ;
        RECT  3.70 0.96 3.86 2.20 ;
        RECT  3.47 1.92 3.86 2.20 ;
        RECT  4.07 0.44 4.35 0.72 ;
        RECT  3.15 0.56 4.35 0.72 ;
        RECT  3.15 0.56 3.31 1.12 ;
        RECT  2.43 0.96 3.31 1.12 ;
        RECT  2.43 0.96 2.71 1.24 ;
        RECT  2.50 0.96 2.66 2.20 ;
        RECT  2.43 1.92 2.71 2.20 ;
        RECT  2.43 2.04 3.31 2.20 ;
        RECT  3.15 2.04 3.31 2.64 ;
        RECT  3.15 2.48 4.25 2.64 ;
        RECT  3.97 2.48 4.25 2.76 ;
        RECT  5.59 0.88 5.91 1.16 ;
        RECT  5.59 0.88 5.75 2.00 ;
        RECT  5.25 1.84 6.23 2.00 ;
        RECT  5.25 1.84 5.53 2.12 ;
        RECT  5.95 1.84 6.23 2.12 ;
        RECT  6.15 0.88 6.43 1.16 ;
        RECT  6.27 0.88 6.43 1.58 ;
        RECT  7.11 1.14 7.39 1.58 ;
        RECT  6.27 1.42 7.39 1.58 ;
        RECT  6.39 1.42 6.55 2.12 ;
        RECT  6.39 1.84 6.75 2.12 ;
        RECT  4.75 0.50 8.15 0.66 ;
        RECT  7.87 0.50 8.15 0.78 ;
        RECT  4.63 0.86 4.91 1.14 ;
        RECT  4.75 0.50 4.91 1.14 ;
        RECT  4.07 0.98 4.91 1.14 ;
        RECT  4.07 0.96 4.35 1.24 ;
        RECT  4.29 0.98 4.45 2.12 ;
        RECT  4.29 1.84 4.57 2.12 ;
        RECT  9.13 0.50 9.41 0.78 ;
        RECT  6.67 0.82 7.71 0.98 ;
        RECT  6.67 0.82 6.95 1.16 ;
        RECT  9.13 0.50 9.29 1.16 ;
        RECT  7.55 1.00 9.29 1.16 ;
        RECT  7.55 0.96 7.91 1.24 ;
        RECT  7.85 1.00 8.01 2.12 ;
        RECT  6.99 1.84 7.27 2.12 ;
        RECT  7.85 1.84 8.19 2.12 ;
        RECT  6.99 1.96 8.19 2.12 ;
        RECT  5.07 0.86 5.43 1.14 ;
        RECT  9.67 0.96 10.11 1.24 ;
        RECT  5.07 0.86 5.23 1.48 ;
        RECT  8.35 1.52 9.83 1.68 ;
        RECT  4.81 1.84 5.09 2.12 ;
        RECT  9.67 0.96 9.83 2.12 ;
        RECT  9.53 1.84 9.83 2.12 ;
        RECT  4.93 1.32 5.09 2.44 ;
        RECT  8.35 1.52 8.51 2.44 ;
        RECT  4.93 2.28 8.51 2.44 ;
        RECT  10.31 0.88 10.73 1.16 ;
        RECT  10.57 1.46 12.11 1.62 ;
        RECT  11.83 1.40 12.11 1.68 ;
        RECT  10.57 0.88 10.73 2.12 ;
        RECT  10.57 1.84 10.85 2.12 ;
        RECT  12.11 0.88 12.47 1.16 ;
        RECT  12.31 0.88 12.47 2.16 ;
        RECT  12.31 1.88 12.59 2.16 ;
        RECT  11.82 2.00 12.59 2.16 ;
        RECT  11.82 2.00 11.98 2.76 ;
        RECT  11.70 2.48 11.98 2.76 ;
    END
END DFFDRSZSP2V1_0

MACRO DFFDRSZSP1V1_0
    CLASS CORE ;
    FOREIGN DFFDRSZSP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 25.99  LAYER ME1  ;
        ANTENNADIFFAREA 10.80  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.60  LAYER ME1  ;
        ANTENNAMAXAREACAR 42.97  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.77 1.89 14.05 2.17 ;
        RECT  13.77 0.88 14.05 1.16 ;
        RECT  13.77 0.88 13.94 2.17 ;
        RECT  13.66 1.46 13.94 1.74 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 25.68  LAYER ME1  ;
        ANTENNADIFFAREA 10.80  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.60  LAYER ME1  ;
        ANTENNAMAXAREACAR 42.46  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.85 1.46 13.14 1.74 ;
        RECT  12.73 1.89 13.01 2.17 ;
        RECT  12.85 0.88 13.01 2.17 ;
        RECT  12.73 0.88 13.01 1.16 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.20  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.83  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.81 1.19 2.25 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  0.91 0.81 1.19 1.09 ;
        END
    END D
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.99 1.40 10.41 1.68 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.24 1.40 3.54 1.76 ;
        END
    END CK
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.66 0.44 11.94 0.94 ;
        RECT  11.45 0.44 11.94 0.72 ;
        END
    END SB
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END SEL
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.87  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 12.90  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.06 1.46 2.34 1.74 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.81 2.23 2.25 ;
        RECT  1.95 0.81 2.23 1.09 ;
        END
    END TD
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 14.40 3.48 ;
        RECT  13.94 2.88 14.22 3.48 ;
        RECT  13.25 1.89 13.53 2.17 ;
        RECT  13.31 1.89 13.47 3.48 ;
        RECT  11.93 2.52 12.21 3.48 ;
        RECT  11.09 1.84 11.37 2.12 ;
        RECT  11.15 1.84 11.31 3.48 ;
        RECT  10.05 1.84 10.33 2.12 ;
        RECT  10.11 1.84 10.27 3.48 ;
        RECT  8.77 1.96 9.29 2.12 ;
        RECT  9.01 1.84 9.29 2.12 ;
        RECT  8.65 2.52 8.93 3.48 ;
        RECT  8.77 1.96 8.93 3.48 ;
        RECT  2.71 2.52 2.99 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 14.40 0.28 ;
        RECT  13.94 -0.28 14.22 0.32 ;
        RECT  13.25 0.88 13.53 1.16 ;
        RECT  13.31 -0.28 13.47 1.16 ;
        RECT  11.08 0.88 11.43 1.16 ;
        RECT  11.08 -0.28 11.24 1.16 ;
        RECT  8.69 -0.28 8.97 0.68 ;
        RECT  2.71 -0.28 2.99 0.68 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  1.55 1.97 1.71 2.57 ;
        RECT  1.55 2.41 2.37 2.57 ;
        RECT  2.09 2.41 2.37 2.69 ;
        RECT  3.47 0.96 3.86 1.24 ;
        RECT  3.70 1.46 4.02 1.74 ;
        RECT  3.70 0.96 3.86 2.20 ;
        RECT  3.47 1.92 3.86 2.20 ;
        RECT  4.07 0.44 4.35 0.72 ;
        RECT  3.15 0.56 4.35 0.72 ;
        RECT  3.15 0.56 3.31 1.12 ;
        RECT  2.43 0.96 3.31 1.12 ;
        RECT  2.43 0.96 2.71 1.24 ;
        RECT  2.50 0.96 2.66 2.20 ;
        RECT  2.43 1.92 2.71 2.20 ;
        RECT  2.43 2.04 3.31 2.20 ;
        RECT  3.15 2.04 3.31 2.64 ;
        RECT  3.15 2.48 4.25 2.64 ;
        RECT  3.97 2.48 4.25 2.76 ;
        RECT  5.59 0.88 5.91 1.16 ;
        RECT  5.59 0.88 5.75 2.00 ;
        RECT  5.25 1.84 6.23 2.00 ;
        RECT  5.25 1.84 5.53 2.12 ;
        RECT  5.95 1.84 6.23 2.12 ;
        RECT  6.15 0.88 6.43 1.16 ;
        RECT  6.27 0.88 6.43 1.58 ;
        RECT  7.11 1.14 7.39 1.58 ;
        RECT  6.27 1.42 7.39 1.58 ;
        RECT  6.39 1.42 6.55 2.12 ;
        RECT  6.39 1.84 6.75 2.12 ;
        RECT  4.75 0.50 8.15 0.66 ;
        RECT  7.87 0.50 8.15 0.78 ;
        RECT  4.63 0.86 4.91 1.14 ;
        RECT  4.75 0.50 4.91 1.14 ;
        RECT  4.07 0.98 4.91 1.14 ;
        RECT  4.07 0.96 4.35 1.24 ;
        RECT  4.29 0.98 4.45 2.12 ;
        RECT  4.29 1.84 4.57 2.12 ;
        RECT  9.13 0.50 9.41 0.78 ;
        RECT  6.67 0.82 7.71 0.98 ;
        RECT  6.67 0.82 6.95 1.16 ;
        RECT  9.13 0.50 9.29 1.16 ;
        RECT  7.55 1.00 9.29 1.16 ;
        RECT  7.55 0.96 7.91 1.24 ;
        RECT  7.85 1.00 8.01 2.12 ;
        RECT  6.99 1.84 7.27 2.12 ;
        RECT  7.85 1.84 8.19 2.12 ;
        RECT  6.99 1.96 8.19 2.12 ;
        RECT  5.07 0.86 5.43 1.14 ;
        RECT  9.67 0.96 10.11 1.24 ;
        RECT  5.07 0.86 5.23 1.48 ;
        RECT  8.35 1.52 9.83 1.68 ;
        RECT  4.81 1.84 5.09 2.12 ;
        RECT  9.67 0.96 9.83 2.12 ;
        RECT  9.53 1.84 9.83 2.12 ;
        RECT  4.93 1.32 5.09 2.44 ;
        RECT  8.35 1.52 8.51 2.44 ;
        RECT  4.93 2.28 8.51 2.44 ;
        RECT  10.31 0.88 10.73 1.16 ;
        RECT  10.57 1.46 12.11 1.62 ;
        RECT  11.83 1.40 12.11 1.68 ;
        RECT  10.57 0.88 10.73 2.12 ;
        RECT  10.57 1.84 10.85 2.12 ;
        RECT  12.11 0.88 12.43 1.16 ;
        RECT  12.27 0.88 12.43 2.16 ;
        RECT  11.93 2.00 12.53 2.16 ;
        RECT  11.93 2.00 12.21 2.28 ;
        RECT  12.37 2.00 12.53 2.64 ;
        RECT  12.37 2.48 12.91 2.64 ;
        RECT  12.63 2.48 12.91 2.76 ;
    END
END DFFDRSZSP1V1_0

MACRO DFFDRSSP8V1_0
    CLASS CORE ;
    FOREIGN DFFDRSSP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 29.68  LAYER ME1  ;
        ANTENNADIFFAREA 15.03  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.56  LAYER ME1  ;
        ANTENNAMAXAREACAR 19.08  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.22 1.88 14.50 2.48 ;
        RECT  14.22 0.64 14.50 1.24 ;
        RECT  14.22 0.64 14.38 2.48 ;
        RECT  13.26 1.52 14.38 1.68 ;
        RECT  13.26 1.46 13.54 1.74 ;
        RECT  13.18 1.88 13.46 2.48 ;
        RECT  13.26 0.64 13.46 2.48 ;
        RECT  13.18 0.64 13.46 1.24 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.40 0.70 1.76 ;
        END
    END D
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.66 1.40 8.08 1.68 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.40 1.16 1.76 ;
        END
    END CK
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.26 0.44 9.54 0.94 ;
        RECT  9.07 0.44 9.54 0.72 ;
        END
    END SB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 29.68  LAYER ME1  ;
        ANTENNADIFFAREA 14.79  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.56  LAYER ME1  ;
        ANTENNAMAXAREACAR 19.08  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.14 1.88 12.42 2.48 ;
        RECT  12.14 0.64 12.42 1.24 ;
        RECT  12.14 0.64 12.30 2.48 ;
        RECT  11.22 1.52 12.30 1.68 ;
        RECT  11.22 1.46 11.54 1.74 ;
        RECT  11.10 1.88 11.38 2.48 ;
        RECT  11.22 0.64 11.38 2.48 ;
        RECT  11.10 0.64 11.38 1.24 ;
        END
    END Q
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 15.20 0.28 ;
        RECT  14.74 0.64 15.02 1.24 ;
        RECT  14.74 -0.28 15.02 0.32 ;
        RECT  14.80 -0.28 14.96 1.24 ;
        RECT  13.70 0.64 13.98 1.24 ;
        RECT  13.76 -0.28 13.92 1.24 ;
        RECT  12.66 0.64 12.94 1.24 ;
        RECT  12.72 -0.28 12.88 1.24 ;
        RECT  11.62 0.64 11.90 1.24 ;
        RECT  11.68 -0.28 11.84 1.24 ;
        RECT  10.58 0.64 10.86 1.24 ;
        RECT  10.64 -0.28 10.80 1.24 ;
        RECT  8.75 0.88 9.10 1.16 ;
        RECT  8.75 -0.28 8.91 1.16 ;
        RECT  6.36 -0.28 6.64 0.68 ;
        RECT  0.38 -0.28 0.66 0.68 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 15.20 3.48 ;
        RECT  14.74 2.88 15.02 3.48 ;
        RECT  14.74 1.88 15.02 2.48 ;
        RECT  14.80 1.88 14.96 3.48 ;
        RECT  13.70 1.88 13.98 2.48 ;
        RECT  13.76 1.88 13.92 3.48 ;
        RECT  12.66 1.88 12.94 2.48 ;
        RECT  12.72 1.88 12.88 3.48 ;
        RECT  11.62 1.88 11.90 2.48 ;
        RECT  11.68 1.88 11.84 3.48 ;
        RECT  10.58 1.88 10.86 2.48 ;
        RECT  10.64 1.88 10.80 3.48 ;
        RECT  9.98 2.40 10.26 3.48 ;
        RECT  8.76 1.84 9.04 2.12 ;
        RECT  8.82 1.84 8.98 3.48 ;
        RECT  7.72 1.84 8.00 2.12 ;
        RECT  7.78 1.84 7.94 3.48 ;
        RECT  6.44 1.96 6.96 2.12 ;
        RECT  6.68 1.84 6.96 2.12 ;
        RECT  6.32 2.52 6.60 3.48 ;
        RECT  6.44 1.96 6.60 3.48 ;
        RECT  0.38 2.48 0.66 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  1.14 0.96 1.48 1.24 ;
        RECT  1.32 1.46 1.64 1.74 ;
        RECT  1.32 0.96 1.48 2.20 ;
        RECT  1.14 1.92 1.48 2.20 ;
        RECT  1.74 0.44 2.02 0.72 ;
        RECT  0.82 0.56 2.02 0.72 ;
        RECT  0.82 0.56 0.98 1.12 ;
        RECT  0.08 0.96 0.98 1.12 ;
        RECT  0.08 0.96 0.38 1.24 ;
        RECT  0.08 0.96 0.24 2.20 ;
        RECT  0.08 1.92 0.38 2.20 ;
        RECT  0.08 2.04 0.98 2.20 ;
        RECT  0.82 2.04 0.98 2.64 ;
        RECT  0.82 2.48 1.92 2.64 ;
        RECT  1.64 2.48 1.92 2.76 ;
        RECT  3.26 0.88 3.58 1.16 ;
        RECT  3.26 0.88 3.42 2.00 ;
        RECT  2.92 1.84 3.90 2.00 ;
        RECT  2.92 1.84 3.20 2.12 ;
        RECT  3.62 1.84 3.90 2.12 ;
        RECT  3.82 0.88 4.10 1.16 ;
        RECT  3.94 0.88 4.10 1.58 ;
        RECT  4.78 1.14 5.06 1.58 ;
        RECT  3.94 1.42 5.06 1.58 ;
        RECT  4.06 1.42 4.22 2.12 ;
        RECT  4.06 1.84 4.42 2.12 ;
        RECT  2.42 0.50 5.82 0.66 ;
        RECT  5.54 0.50 5.82 0.78 ;
        RECT  2.30 0.86 2.58 1.14 ;
        RECT  2.42 0.50 2.58 1.14 ;
        RECT  1.74 0.98 2.58 1.14 ;
        RECT  1.74 0.96 2.02 1.24 ;
        RECT  1.96 0.98 2.12 2.12 ;
        RECT  1.96 1.84 2.24 2.12 ;
        RECT  6.80 0.50 7.08 0.78 ;
        RECT  4.34 0.82 5.38 0.98 ;
        RECT  4.34 0.82 4.62 1.16 ;
        RECT  6.80 0.50 6.96 1.16 ;
        RECT  5.22 1.00 6.96 1.16 ;
        RECT  5.22 0.96 5.58 1.24 ;
        RECT  5.52 1.00 5.68 2.12 ;
        RECT  4.66 1.84 4.94 2.12 ;
        RECT  5.52 1.84 5.86 2.12 ;
        RECT  4.66 1.96 5.86 2.12 ;
        RECT  2.74 0.86 3.10 1.14 ;
        RECT  7.34 0.96 7.78 1.24 ;
        RECT  2.74 0.86 2.90 1.48 ;
        RECT  6.02 1.52 7.50 1.68 ;
        RECT  2.48 1.84 2.76 2.12 ;
        RECT  7.34 0.96 7.50 2.12 ;
        RECT  7.20 1.84 7.50 2.12 ;
        RECT  2.60 1.32 2.76 2.44 ;
        RECT  6.02 1.52 6.18 2.44 ;
        RECT  2.60 2.28 6.18 2.44 ;
        RECT  7.98 0.88 8.40 1.16 ;
        RECT  8.24 1.46 9.78 1.62 ;
        RECT  9.50 1.40 9.78 1.68 ;
        RECT  8.24 0.88 8.40 2.12 ;
        RECT  8.24 1.84 8.52 2.12 ;
        RECT  9.78 0.88 10.14 1.16 ;
        RECT  9.98 0.88 10.14 2.16 ;
        RECT  9.49 1.96 10.26 2.12 ;
        RECT  9.98 1.88 10.26 2.16 ;
        RECT  9.49 1.96 9.65 2.76 ;
        RECT  9.37 2.48 9.65 2.76 ;
    END
END DFFDRSSP8V1_0

MACRO DFFDRSSP4V1_0
    CLASS CORE ;
    FOREIGN DFFDRSSP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 13.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 25.43  LAYER ME1  ;
        ANTENNADIFFAREA 11.99  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.98  LAYER ME1  ;
        ANTENNAMAXAREACAR 25.97  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.14 1.88 12.42 2.48 ;
        RECT  12.14 0.64 12.42 1.24 ;
        RECT  12.14 0.64 12.34 2.48 ;
        RECT  12.06 1.46 12.34 1.74 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 25.43  LAYER ME1  ;
        ANTENNADIFFAREA 11.75  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.98  LAYER ME1  ;
        ANTENNAMAXAREACAR 25.97  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.22 1.46 11.54 1.74 ;
        RECT  11.10 1.88 11.38 2.48 ;
        RECT  11.22 0.64 11.38 2.48 ;
        RECT  11.10 0.64 11.38 1.24 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.26 0.44 9.54 0.94 ;
        RECT  9.07 0.44 9.54 0.72 ;
        END
    END SB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.40 1.16 1.76 ;
        END
    END CK
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.66 1.40 8.08 1.68 ;
        END
    END RB
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.40 0.70 1.76 ;
        END
    END D
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 13.20 0.28 ;
        RECT  12.72 -0.28 13.02 0.32 ;
        RECT  12.66 0.64 12.94 1.24 ;
        RECT  12.72 -0.28 12.88 1.24 ;
        RECT  11.62 0.64 11.90 1.24 ;
        RECT  11.68 -0.28 11.84 1.24 ;
        RECT  10.58 0.64 10.86 1.24 ;
        RECT  10.64 -0.28 10.80 1.24 ;
        RECT  8.75 0.88 9.10 1.16 ;
        RECT  8.75 -0.28 8.91 1.16 ;
        RECT  6.36 -0.28 6.64 0.68 ;
        RECT  0.38 -0.28 0.66 0.68 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 13.20 3.48 ;
        RECT  12.72 2.88 13.02 3.48 ;
        RECT  12.66 1.88 12.94 2.48 ;
        RECT  12.72 1.88 12.88 3.48 ;
        RECT  11.62 1.88 11.90 2.48 ;
        RECT  11.68 1.88 11.84 3.48 ;
        RECT  10.58 1.88 10.86 2.48 ;
        RECT  10.64 1.88 10.80 3.48 ;
        RECT  9.98 2.40 10.26 3.48 ;
        RECT  8.76 1.84 9.04 2.12 ;
        RECT  8.82 1.84 8.98 3.48 ;
        RECT  7.72 1.84 8.00 2.12 ;
        RECT  7.78 1.84 7.94 3.48 ;
        RECT  6.44 1.96 6.96 2.12 ;
        RECT  6.68 1.84 6.96 2.12 ;
        RECT  6.32 2.52 6.60 3.48 ;
        RECT  6.44 1.96 6.60 3.48 ;
        RECT  0.38 2.48 0.66 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  1.14 0.96 1.48 1.24 ;
        RECT  1.32 1.46 1.64 1.74 ;
        RECT  1.32 0.96 1.48 2.20 ;
        RECT  1.14 1.92 1.48 2.20 ;
        RECT  1.74 0.44 2.02 0.72 ;
        RECT  0.82 0.56 2.02 0.72 ;
        RECT  0.82 0.56 0.98 1.12 ;
        RECT  0.08 0.96 0.98 1.12 ;
        RECT  0.08 0.96 0.38 1.24 ;
        RECT  0.08 0.96 0.24 2.20 ;
        RECT  0.08 1.92 0.38 2.20 ;
        RECT  0.08 2.04 0.98 2.20 ;
        RECT  0.82 2.04 0.98 2.64 ;
        RECT  0.82 2.48 1.92 2.64 ;
        RECT  1.64 2.48 1.92 2.76 ;
        RECT  3.26 0.88 3.58 1.16 ;
        RECT  3.26 0.88 3.42 2.00 ;
        RECT  2.92 1.84 3.90 2.00 ;
        RECT  2.92 1.84 3.20 2.12 ;
        RECT  3.62 1.84 3.90 2.12 ;
        RECT  3.82 0.88 4.10 1.16 ;
        RECT  3.94 0.88 4.10 1.58 ;
        RECT  4.78 1.14 5.06 1.58 ;
        RECT  3.94 1.42 5.06 1.58 ;
        RECT  4.06 1.42 4.22 2.12 ;
        RECT  4.06 1.84 4.42 2.12 ;
        RECT  2.42 0.50 5.82 0.66 ;
        RECT  5.54 0.50 5.82 0.78 ;
        RECT  2.30 0.86 2.58 1.14 ;
        RECT  2.42 0.50 2.58 1.14 ;
        RECT  1.74 0.98 2.58 1.14 ;
        RECT  1.74 0.96 2.02 1.24 ;
        RECT  1.96 0.98 2.12 2.12 ;
        RECT  1.96 1.84 2.24 2.12 ;
        RECT  6.80 0.50 7.08 0.78 ;
        RECT  4.34 0.82 5.38 0.98 ;
        RECT  4.34 0.82 4.62 1.16 ;
        RECT  6.80 0.50 6.96 1.16 ;
        RECT  5.22 1.00 6.96 1.16 ;
        RECT  5.22 0.96 5.58 1.24 ;
        RECT  5.52 1.00 5.68 2.12 ;
        RECT  4.66 1.84 4.94 2.12 ;
        RECT  5.52 1.84 5.86 2.12 ;
        RECT  4.66 1.96 5.86 2.12 ;
        RECT  2.74 0.86 3.10 1.14 ;
        RECT  7.34 0.96 7.78 1.24 ;
        RECT  2.74 0.86 2.90 1.48 ;
        RECT  6.02 1.52 7.50 1.68 ;
        RECT  2.48 1.84 2.76 2.12 ;
        RECT  7.34 0.96 7.50 2.12 ;
        RECT  7.20 1.84 7.50 2.12 ;
        RECT  2.60 1.32 2.76 2.44 ;
        RECT  6.02 1.52 6.18 2.44 ;
        RECT  2.60 2.28 6.18 2.44 ;
        RECT  7.98 0.88 8.40 1.16 ;
        RECT  8.24 1.46 9.78 1.62 ;
        RECT  9.50 1.40 9.78 1.68 ;
        RECT  8.24 0.88 8.40 2.12 ;
        RECT  8.24 1.84 8.52 2.12 ;
        RECT  9.78 0.88 10.14 1.16 ;
        RECT  9.98 0.88 10.14 2.16 ;
        RECT  9.49 1.96 10.26 2.12 ;
        RECT  9.98 1.88 10.26 2.16 ;
        RECT  9.49 1.96 9.65 2.76 ;
        RECT  9.37 2.48 9.65 2.76 ;
    END
END DFFDRSSP4V1_0

MACRO DFFDRSSP2V1_0
    CLASS CORE ;
    FOREIGN DFFDRSSP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 23.16  LAYER ME1  ;
        ANTENNADIFFAREA 10.40  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.69  LAYER ME1  ;
        ANTENNAMAXAREACAR 33.50  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.66 1.46 11.92 1.74 ;
        RECT  11.62 1.84 11.90 2.44 ;
        RECT  11.66 0.64 11.90 2.44 ;
        RECT  11.62 0.64 11.90 1.24 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 23.16  LAYER ME1  ;
        ANTENNADIFFAREA 10.40  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.69  LAYER ME1  ;
        ANTENNAMAXAREACAR 33.50  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.58 1.84 10.86 2.44 ;
        RECT  10.58 0.64 10.86 1.24 ;
        RECT  10.58 0.64 10.74 2.44 ;
        RECT  10.46 1.46 10.74 1.74 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.40 0.70 1.76 ;
        END
    END D
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.66 1.40 8.08 1.68 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.40 1.16 1.76 ;
        END
    END CK
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.26 0.44 9.54 0.94 ;
        RECT  9.07 0.44 9.54 0.72 ;
        END
    END SB
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 12.00 3.48 ;
        RECT  11.54 2.88 11.82 3.48 ;
        RECT  11.10 1.84 11.38 2.44 ;
        RECT  11.16 1.84 11.32 3.48 ;
        RECT  9.98 2.40 10.26 3.48 ;
        RECT  8.76 1.84 9.04 2.12 ;
        RECT  8.82 1.84 8.98 3.48 ;
        RECT  7.72 1.84 8.00 2.12 ;
        RECT  7.78 1.84 7.94 3.48 ;
        RECT  6.44 1.96 6.96 2.12 ;
        RECT  6.68 1.84 6.96 2.12 ;
        RECT  6.32 2.52 6.60 3.48 ;
        RECT  6.44 1.96 6.60 3.48 ;
        RECT  0.38 2.48 0.66 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 12.00 0.28 ;
        RECT  11.54 -0.28 11.82 0.32 ;
        RECT  11.10 0.64 11.38 1.24 ;
        RECT  11.16 -0.28 11.32 1.24 ;
        RECT  8.75 0.88 9.10 1.16 ;
        RECT  8.75 -0.28 8.91 1.16 ;
        RECT  6.36 -0.28 6.64 0.68 ;
        RECT  0.38 -0.28 0.66 0.68 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  1.14 0.96 1.48 1.24 ;
        RECT  1.32 1.46 1.64 1.74 ;
        RECT  1.32 0.96 1.48 2.20 ;
        RECT  1.14 1.92 1.48 2.20 ;
        RECT  1.74 0.44 2.02 0.72 ;
        RECT  0.82 0.56 2.02 0.72 ;
        RECT  0.82 0.56 0.98 1.12 ;
        RECT  0.08 0.96 0.98 1.12 ;
        RECT  0.08 0.96 0.38 1.24 ;
        RECT  0.08 0.96 0.24 2.20 ;
        RECT  0.08 1.92 0.38 2.20 ;
        RECT  0.08 2.04 0.98 2.20 ;
        RECT  0.82 2.04 0.98 2.64 ;
        RECT  0.82 2.48 1.92 2.64 ;
        RECT  1.64 2.48 1.92 2.76 ;
        RECT  3.26 0.88 3.58 1.16 ;
        RECT  3.26 0.88 3.42 2.00 ;
        RECT  2.92 1.84 3.90 2.00 ;
        RECT  2.92 1.84 3.20 2.12 ;
        RECT  3.62 1.84 3.90 2.12 ;
        RECT  3.82 0.88 4.10 1.16 ;
        RECT  3.94 0.88 4.10 1.58 ;
        RECT  4.78 1.14 5.06 1.58 ;
        RECT  3.94 1.42 5.06 1.58 ;
        RECT  4.06 1.42 4.22 2.12 ;
        RECT  4.06 1.84 4.42 2.12 ;
        RECT  2.42 0.50 5.82 0.66 ;
        RECT  5.54 0.50 5.82 0.78 ;
        RECT  2.30 0.86 2.58 1.14 ;
        RECT  2.42 0.50 2.58 1.14 ;
        RECT  1.74 0.98 2.58 1.14 ;
        RECT  1.74 0.96 2.02 1.24 ;
        RECT  1.96 0.98 2.12 2.12 ;
        RECT  1.96 1.84 2.24 2.12 ;
        RECT  6.80 0.50 7.08 0.78 ;
        RECT  4.34 0.82 5.38 0.98 ;
        RECT  4.34 0.82 4.62 1.16 ;
        RECT  6.80 0.50 6.96 1.16 ;
        RECT  5.22 1.00 6.96 1.16 ;
        RECT  5.22 0.96 5.58 1.24 ;
        RECT  5.52 1.00 5.68 2.12 ;
        RECT  4.66 1.84 4.94 2.12 ;
        RECT  5.52 1.84 5.86 2.12 ;
        RECT  4.66 1.96 5.86 2.12 ;
        RECT  2.74 0.86 3.10 1.14 ;
        RECT  7.34 0.96 7.78 1.24 ;
        RECT  2.74 0.86 2.90 1.48 ;
        RECT  6.02 1.52 7.50 1.68 ;
        RECT  2.48 1.84 2.76 2.12 ;
        RECT  7.34 0.96 7.50 2.12 ;
        RECT  7.20 1.84 7.50 2.12 ;
        RECT  2.60 1.32 2.76 2.44 ;
        RECT  6.02 1.52 6.18 2.44 ;
        RECT  2.60 2.28 6.18 2.44 ;
        RECT  7.98 0.88 8.40 1.16 ;
        RECT  8.24 1.46 9.78 1.62 ;
        RECT  9.50 1.40 9.78 1.68 ;
        RECT  8.24 0.88 8.40 2.12 ;
        RECT  8.24 1.84 8.52 2.12 ;
        RECT  9.78 0.88 10.14 1.16 ;
        RECT  9.98 0.88 10.14 2.16 ;
        RECT  9.49 1.96 10.26 2.12 ;
        RECT  9.98 1.88 10.26 2.16 ;
        RECT  9.49 1.96 9.65 2.76 ;
        RECT  9.37 2.48 9.65 2.76 ;
    END
END DFFDRSSP2V1_0

MACRO DFFDRSSP1V1_0
    CLASS CORE ;
    FOREIGN DFFDRSSP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.26 0.44 9.54 0.94 ;
        RECT  9.07 0.44 9.54 0.72 ;
        END
    END SB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 22.70  LAYER ME1  ;
        ANTENNADIFFAREA 9.64  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.54  LAYER ME1  ;
        ANTENNAMAXAREACAR 42.23  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.46 1.46 10.74 1.74 ;
        RECT  10.36 1.84 10.64 2.12 ;
        RECT  10.46 0.88 10.64 2.12 ;
        RECT  10.36 0.88 10.64 1.16 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 22.40  LAYER ME1  ;
        ANTENNADIFFAREA 9.64  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.54  LAYER ME1  ;
        ANTENNAMAXAREACAR 41.67  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.40 1.84 11.68 2.12 ;
        RECT  11.40 0.88 11.68 1.16 ;
        RECT  11.40 0.88 11.56 2.12 ;
        RECT  11.29 1.46 11.56 1.74 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.40 0.70 1.76 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.40 1.16 1.76 ;
        END
    END CK
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.66 1.40 8.08 1.68 ;
        END
    END RB
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 12.00 0.28 ;
        RECT  11.54 -0.28 11.82 0.32 ;
        RECT  10.88 0.88 11.16 1.16 ;
        RECT  10.94 -0.28 11.10 1.16 ;
        RECT  8.75 0.88 9.10 1.16 ;
        RECT  8.75 -0.28 8.91 1.16 ;
        RECT  6.36 -0.28 6.64 0.68 ;
        RECT  0.38 -0.28 0.66 0.68 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 12.00 3.48 ;
        RECT  11.54 2.88 11.82 3.48 ;
        RECT  10.88 1.84 11.16 2.12 ;
        RECT  10.94 1.84 11.10 3.48 ;
        RECT  9.60 2.52 9.88 3.48 ;
        RECT  8.76 1.84 9.04 2.12 ;
        RECT  8.82 1.84 8.98 3.48 ;
        RECT  7.72 1.84 8.00 2.12 ;
        RECT  7.78 1.84 7.94 3.48 ;
        RECT  6.44 1.96 6.96 2.12 ;
        RECT  6.68 1.84 6.96 2.12 ;
        RECT  6.32 2.52 6.60 3.48 ;
        RECT  6.44 1.96 6.60 3.48 ;
        RECT  0.38 2.48 0.66 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  1.14 0.96 1.48 1.24 ;
        RECT  1.32 1.46 1.64 1.74 ;
        RECT  1.32 0.96 1.48 2.20 ;
        RECT  1.14 1.92 1.48 2.20 ;
        RECT  1.74 0.44 2.02 0.72 ;
        RECT  0.82 0.56 2.02 0.72 ;
        RECT  0.82 0.56 0.98 1.12 ;
        RECT  0.08 0.96 0.98 1.12 ;
        RECT  0.08 0.96 0.38 1.24 ;
        RECT  0.08 0.96 0.24 2.20 ;
        RECT  0.08 1.92 0.38 2.20 ;
        RECT  0.08 2.04 0.98 2.20 ;
        RECT  0.82 2.04 0.98 2.64 ;
        RECT  0.82 2.48 1.92 2.64 ;
        RECT  1.64 2.48 1.92 2.76 ;
        RECT  3.26 0.88 3.58 1.16 ;
        RECT  3.26 0.88 3.42 2.00 ;
        RECT  2.92 1.84 3.90 2.00 ;
        RECT  2.92 1.84 3.20 2.12 ;
        RECT  3.62 1.84 3.90 2.12 ;
        RECT  3.82 0.88 4.10 1.16 ;
        RECT  3.94 0.88 4.10 1.58 ;
        RECT  4.78 1.14 5.06 1.58 ;
        RECT  3.94 1.42 5.06 1.58 ;
        RECT  4.06 1.42 4.22 2.12 ;
        RECT  4.06 1.84 4.42 2.12 ;
        RECT  2.42 0.50 5.82 0.66 ;
        RECT  5.54 0.50 5.82 0.78 ;
        RECT  2.30 0.86 2.58 1.14 ;
        RECT  2.42 0.50 2.58 1.14 ;
        RECT  1.74 0.98 2.58 1.14 ;
        RECT  1.74 0.96 2.02 1.24 ;
        RECT  1.96 0.98 2.12 2.12 ;
        RECT  1.96 1.84 2.24 2.12 ;
        RECT  6.80 0.50 7.08 0.78 ;
        RECT  4.34 0.82 5.38 0.98 ;
        RECT  4.34 0.82 4.62 1.16 ;
        RECT  6.80 0.50 6.96 1.16 ;
        RECT  5.22 1.00 6.96 1.16 ;
        RECT  5.22 0.96 5.58 1.24 ;
        RECT  5.52 1.00 5.68 2.12 ;
        RECT  4.66 1.84 4.94 2.12 ;
        RECT  5.52 1.84 5.86 2.12 ;
        RECT  4.66 1.96 5.86 2.12 ;
        RECT  2.74 0.86 3.10 1.14 ;
        RECT  7.34 0.96 7.78 1.24 ;
        RECT  2.74 0.86 2.90 1.48 ;
        RECT  6.02 1.52 7.50 1.68 ;
        RECT  2.48 1.84 2.76 2.12 ;
        RECT  7.34 0.96 7.50 2.12 ;
        RECT  7.20 1.84 7.50 2.12 ;
        RECT  2.60 1.32 2.76 2.44 ;
        RECT  6.02 1.52 6.18 2.44 ;
        RECT  2.60 2.28 6.18 2.44 ;
        RECT  7.98 0.88 8.40 1.16 ;
        RECT  8.24 1.46 9.78 1.62 ;
        RECT  9.50 1.40 9.78 1.68 ;
        RECT  8.24 0.88 8.40 2.12 ;
        RECT  8.24 1.84 8.52 2.12 ;
        RECT  9.78 0.88 10.10 1.16 ;
        RECT  9.94 0.88 10.10 2.16 ;
        RECT  9.60 2.00 10.20 2.16 ;
        RECT  9.60 2.00 9.88 2.28 ;
        RECT  10.04 2.00 10.20 2.64 ;
        RECT  10.04 2.48 10.58 2.64 ;
        RECT  10.30 2.48 10.58 2.76 ;
    END
END DFFDRSSP1V1_0

MACRO DFFDRSP8V1_1
    CLASS CORE ;
    FOREIGN DFFDRSP8V1_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 13.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 27.03  LAYER ME1  ;
        ANTENNADIFFAREA 13.66  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.56  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.38  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.58 1.90 12.86 2.50 ;
        RECT  12.58 0.64 12.86 1.24 ;
        RECT  12.58 0.64 12.74 2.50 ;
        RECT  11.66 1.52 12.74 1.68 ;
        RECT  11.66 1.46 11.94 1.74 ;
        RECT  11.54 1.90 11.82 2.50 ;
        RECT  11.66 0.64 11.82 2.50 ;
        RECT  11.54 0.64 11.82 1.24 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 27.03  LAYER ME1  ;
        ANTENNADIFFAREA 13.40  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.56  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.38  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.50 1.90 10.78 2.50 ;
        RECT  10.50 0.64 10.78 1.24 ;
        RECT  10.50 0.64 10.66 2.50 ;
        RECT  9.58 1.52 10.66 1.68 ;
        RECT  9.58 1.46 9.94 1.74 ;
        RECT  9.46 1.90 9.74 2.50 ;
        RECT  9.58 0.64 9.74 2.50 ;
        RECT  9.46 0.64 9.74 1.24 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.40 0.72 1.76 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.88 1.40 1.20 1.76 ;
        END
    END CK
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.42 2.28 6.80 2.56 ;
        END
    END RB
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 13.60 0.28 ;
        RECT  13.14 -0.28 13.42 0.32 ;
        RECT  13.10 0.64 13.38 1.24 ;
        RECT  13.16 -0.28 13.32 1.24 ;
        RECT  12.06 0.64 12.34 1.24 ;
        RECT  12.12 -0.28 12.28 1.24 ;
        RECT  11.02 0.64 11.30 1.24 ;
        RECT  11.08 -0.28 11.24 1.24 ;
        RECT  9.98 0.64 10.26 1.24 ;
        RECT  10.04 -0.28 10.20 1.24 ;
        RECT  8.94 0.64 9.22 1.24 ;
        RECT  9.00 -0.28 9.16 1.24 ;
        RECT  7.94 0.88 8.22 1.16 ;
        RECT  8.00 -0.28 8.16 1.16 ;
        RECT  4.96 -0.28 5.24 0.72 ;
        RECT  0.38 -0.28 0.66 0.68 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 13.60 3.48 ;
        RECT  13.14 2.88 13.42 3.48 ;
        RECT  13.10 1.90 13.38 2.50 ;
        RECT  13.16 1.90 13.32 3.48 ;
        RECT  12.06 1.90 12.34 2.50 ;
        RECT  12.12 1.90 12.28 3.48 ;
        RECT  11.02 1.90 11.30 2.50 ;
        RECT  11.08 1.90 11.24 3.48 ;
        RECT  9.98 1.90 10.26 2.50 ;
        RECT  10.04 1.90 10.20 3.48 ;
        RECT  8.94 1.90 9.22 2.50 ;
        RECT  9.00 1.90 9.16 3.48 ;
        RECT  7.94 1.84 8.22 2.12 ;
        RECT  8.00 1.84 8.16 3.48 ;
        RECT  7.10 1.84 7.26 3.48 ;
        RECT  6.90 1.84 7.26 2.12 ;
        RECT  6.06 1.84 6.22 3.48 ;
        RECT  5.86 1.84 6.22 2.12 ;
        RECT  0.38 2.48 0.66 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  1.14 0.96 1.52 1.24 ;
        RECT  1.36 1.46 1.64 1.74 ;
        RECT  1.36 0.96 1.52 2.20 ;
        RECT  1.14 1.92 1.52 2.20 ;
        RECT  1.74 0.44 2.02 0.72 ;
        RECT  0.82 0.56 2.02 0.72 ;
        RECT  0.82 0.56 0.98 1.12 ;
        RECT  0.08 0.96 0.98 1.12 ;
        RECT  0.08 0.96 0.38 1.24 ;
        RECT  0.08 0.96 0.24 2.20 ;
        RECT  0.08 1.92 0.38 2.20 ;
        RECT  0.08 2.04 0.98 2.20 ;
        RECT  0.82 2.04 0.98 2.64 ;
        RECT  0.82 2.48 2.02 2.64 ;
        RECT  1.74 2.48 2.02 2.76 ;
        RECT  3.34 0.88 3.62 1.16 ;
        RECT  3.34 0.88 3.50 2.12 ;
        RECT  3.12 1.84 3.50 2.12 ;
        RECT  3.82 1.84 4.10 2.12 ;
        RECT  3.12 1.96 4.10 2.12 ;
        RECT  4.52 0.44 4.80 0.72 ;
        RECT  3.98 0.56 4.80 0.72 ;
        RECT  3.86 0.88 4.14 1.16 ;
        RECT  3.98 0.56 4.14 1.68 ;
        RECT  3.98 1.52 4.42 1.68 ;
        RECT  4.26 1.52 4.42 2.12 ;
        RECT  4.26 1.84 4.62 2.12 ;
        RECT  2.30 0.87 2.58 1.15 ;
        RECT  1.74 0.99 2.58 1.15 ;
        RECT  1.74 0.96 2.02 1.24 ;
        RECT  1.86 0.96 2.02 2.12 ;
        RECT  1.86 1.84 2.14 2.12 ;
        RECT  1.86 1.96 2.44 2.12 ;
        RECT  2.28 1.96 2.44 2.76 ;
        RECT  5.62 2.42 5.90 2.76 ;
        RECT  2.28 2.60 5.90 2.76 ;
        RECT  5.82 0.50 6.10 0.78 ;
        RECT  4.38 0.88 4.66 1.20 ;
        RECT  5.00 0.92 5.28 1.20 ;
        RECT  5.82 0.50 5.98 1.20 ;
        RECT  4.38 1.04 5.98 1.20 ;
        RECT  4.78 1.04 4.94 2.12 ;
        RECT  4.78 1.84 5.14 2.12 ;
        RECT  2.80 0.87 3.10 1.15 ;
        RECT  6.48 0.92 6.76 1.20 ;
        RECT  5.30 1.52 6.64 1.68 ;
        RECT  6.48 0.92 6.64 2.12 ;
        RECT  2.68 1.84 2.96 2.12 ;
        RECT  6.38 1.84 6.66 2.12 ;
        RECT  2.80 0.87 2.96 2.44 ;
        RECT  5.30 1.52 5.46 2.44 ;
        RECT  2.80 2.28 5.46 2.44 ;
        RECT  7.04 0.88 7.32 1.16 ;
        RECT  7.04 1.00 7.58 1.16 ;
        RECT  7.42 1.46 8.42 1.62 ;
        RECT  8.14 1.40 8.42 1.68 ;
        RECT  7.42 1.00 7.58 2.12 ;
        RECT  7.42 1.84 7.70 2.12 ;
        RECT  8.46 0.88 8.74 1.16 ;
        RECT  8.46 1.84 8.74 2.12 ;
        RECT  8.58 0.88 8.74 2.76 ;
        RECT  8.49 2.48 8.77 2.76 ;
    END
END DFFDRSP8V1_1

MACRO DFFDRSP8V1_0
    CLASS CORE ;
    FOREIGN DFFDRSP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 27.31  LAYER ME1  ;
        ANTENNADIFFAREA 12.74  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.79  LAYER ME1  ;
        ANTENNAMAXAREACAR 15.25  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.91 1.92 13.19 2.52 ;
        RECT  12.91 0.64 13.19 1.24 ;
        RECT  12.92 0.64 13.08 2.52 ;
        RECT  11.99 1.52 13.08 1.68 ;
        RECT  11.87 1.92 12.15 2.52 ;
        RECT  11.99 0.64 12.15 2.52 ;
        RECT  11.87 0.64 12.15 1.24 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 27.31  LAYER ME1  ;
        ANTENNADIFFAREA 13.10  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.79  LAYER ME1  ;
        ANTENNAMAXAREACAR 15.25  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.83 1.92 11.11 2.52 ;
        RECT  10.83 0.64 11.11 1.24 ;
        RECT  10.83 0.64 10.99 2.52 ;
        RECT  9.72 1.52 10.99 1.68 ;
        RECT  9.72 1.92 10.07 2.52 ;
        RECT  9.72 0.64 10.07 1.24 ;
        RECT  9.72 0.64 9.88 2.52 ;
        END
    END Q
    PIN RB
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.42  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        ANTENNAMAXAREACAR 3.16  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.71 1.46 9.14 1.74 ;
        RECT  4.62 2.54 6.82 2.70 ;
        RECT  6.54 2.42 6.82 2.70 ;
        RECT  4.62 2.40 4.90 2.70 ;
        END
    END RB
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.66 1.34 1.94 1.76 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.46 1.39 0.74 1.81 ;
        END
    END CK
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 14.00 0.28 ;
        RECT  13.49 -0.28 13.82 0.32 ;
        RECT  13.43 0.64 13.71 1.24 ;
        RECT  13.49 -0.28 13.65 1.24 ;
        RECT  12.39 0.64 12.67 1.24 ;
        RECT  12.45 -0.28 12.61 1.24 ;
        RECT  11.35 0.64 11.63 1.24 ;
        RECT  11.41 -0.28 11.57 1.24 ;
        RECT  10.31 0.64 10.59 1.24 ;
        RECT  10.37 -0.28 10.53 1.24 ;
        RECT  9.27 0.64 9.55 1.24 ;
        RECT  9.33 -0.28 9.49 1.24 ;
        RECT  7.75 0.96 8.03 1.24 ;
        RECT  7.82 -0.28 7.98 1.24 ;
        RECT  4.29 0.76 4.57 1.04 ;
        RECT  4.35 -0.28 4.51 1.04 ;
        RECT  1.64 0.76 1.92 1.04 ;
        RECT  1.70 -0.28 1.86 1.04 ;
        RECT  0.62 0.50 0.90 0.78 ;
        RECT  0.68 -0.28 0.84 0.78 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 14.00 3.48 ;
        RECT  13.49 2.88 13.82 3.48 ;
        RECT  13.43 1.92 13.71 2.52 ;
        RECT  13.49 1.92 13.65 3.48 ;
        RECT  12.39 1.92 12.67 2.52 ;
        RECT  12.45 1.92 12.61 3.48 ;
        RECT  11.35 1.92 11.63 2.52 ;
        RECT  11.41 1.92 11.57 3.48 ;
        RECT  10.31 1.92 10.59 2.52 ;
        RECT  10.38 1.92 10.54 3.48 ;
        RECT  9.27 1.92 9.55 2.52 ;
        RECT  9.33 1.92 9.49 3.48 ;
        RECT  8.77 1.90 9.05 2.18 ;
        RECT  8.83 1.90 8.99 3.48 ;
        RECT  7.73 1.90 8.01 2.18 ;
        RECT  7.79 1.90 7.95 3.48 ;
        RECT  3.76 2.08 5.08 2.24 ;
        RECT  4.80 1.96 5.08 2.24 ;
        RECT  4.30 2.08 4.46 3.48 ;
        RECT  3.76 1.96 4.04 2.24 ;
        RECT  1.64 1.92 1.92 2.20 ;
        RECT  1.72 1.92 1.88 3.48 ;
        RECT  0.62 1.97 0.90 2.25 ;
        RECT  0.68 1.97 0.84 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.07 0.50 0.38 0.78 ;
        RECT  0.07 0.94 1.16 1.10 ;
        RECT  0.88 0.94 1.16 1.22 ;
        RECT  0.07 0.50 0.23 2.25 ;
        RECT  0.07 1.97 0.38 2.25 ;
        RECT  1.14 0.50 1.48 0.78 ;
        RECT  1.14 1.97 1.48 2.25 ;
        RECT  1.32 0.50 1.48 2.70 ;
        RECT  1.28 2.42 1.56 2.70 ;
        RECT  2.16 0.76 2.44 1.04 ;
        RECT  2.22 0.76 2.38 2.20 ;
        RECT  2.16 1.92 2.44 2.20 ;
        RECT  3.20 0.76 3.48 1.04 ;
        RECT  3.26 0.76 3.42 2.20 ;
        RECT  3.20 1.92 3.48 2.20 ;
        RECT  3.32 1.92 3.48 2.62 ;
        RECT  3.32 2.46 4.00 2.62 ;
        RECT  3.72 2.46 4.00 2.74 ;
        RECT  2.80 0.44 3.94 0.60 ;
        RECT  2.80 0.44 2.96 1.04 ;
        RECT  2.68 0.76 2.96 1.04 ;
        RECT  3.78 0.44 3.94 1.36 ;
        RECT  3.78 1.20 5.08 1.36 ;
        RECT  4.80 1.20 5.08 1.48 ;
        RECT  2.74 0.76 2.90 2.20 ;
        RECT  2.68 1.92 2.96 2.20 ;
        RECT  5.04 0.76 5.40 1.04 ;
        RECT  3.59 1.52 3.87 1.80 ;
        RECT  3.59 1.64 5.40 1.80 ;
        RECT  5.24 0.76 5.40 2.24 ;
        RECT  5.24 1.96 5.60 2.24 ;
        RECT  5.76 0.44 7.37 0.60 ;
        RECT  7.09 0.44 7.37 0.72 ;
        RECT  5.56 0.76 5.92 1.04 ;
        RECT  5.76 0.44 5.92 2.24 ;
        RECT  5.76 1.96 6.12 2.24 ;
        RECT  6.69 1.90 6.97 2.24 ;
        RECT  5.76 2.08 6.97 2.24 ;
        RECT  6.08 0.76 6.36 1.12 ;
        RECT  6.08 0.96 7.51 1.12 ;
        RECT  7.21 0.96 7.51 1.24 ;
        RECT  6.21 0.96 6.37 1.81 ;
        RECT  6.21 1.53 6.49 1.81 ;
        RECT  7.21 0.96 7.37 2.18 ;
        RECT  7.21 1.90 7.49 2.18 ;
        RECT  8.79 0.44 9.07 0.72 ;
        RECT  8.33 0.96 8.95 1.12 ;
        RECT  8.79 0.44 8.95 1.24 ;
        RECT  8.65 0.96 8.95 1.24 ;
        RECT  7.55 1.52 8.49 1.68 ;
        RECT  7.55 1.46 7.83 1.74 ;
        RECT  8.33 0.96 8.49 2.18 ;
        RECT  8.25 1.90 8.53 2.18 ;
    END
END DFFDRSP8V1_0

MACRO DFFDRSP4V1_1
    CLASS CORE ;
    FOREIGN DFFDRSP4V1_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.42 2.28 6.80 2.56 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.88 1.40 1.20 1.76 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.40 0.72 1.76 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 22.83  LAYER ME1  ;
        ANTENNADIFFAREA 10.36  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.98  LAYER ME1  ;
        ANTENNAMAXAREACAR 23.31  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.58 1.46 9.94 1.74 ;
        RECT  9.46 1.90 9.74 2.50 ;
        RECT  9.58 0.64 9.74 2.50 ;
        RECT  9.46 0.64 9.74 1.24 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 22.83  LAYER ME1  ;
        ANTENNADIFFAREA 10.62  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.98  LAYER ME1  ;
        ANTENNAMAXAREACAR 23.31  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.50 1.90 10.78 2.50 ;
        RECT  10.50 0.64 10.78 1.24 ;
        RECT  10.50 0.64 10.74 2.50 ;
        RECT  10.46 1.46 10.74 1.74 ;
        END
    END QB
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 11.60 3.48 ;
        RECT  11.08 2.88 11.42 3.48 ;
        RECT  11.02 1.90 11.30 2.50 ;
        RECT  11.08 1.90 11.24 3.48 ;
        RECT  9.98 1.90 10.26 2.50 ;
        RECT  10.04 1.90 10.20 3.48 ;
        RECT  8.94 1.90 9.22 2.50 ;
        RECT  9.00 1.90 9.16 3.48 ;
        RECT  7.94 1.84 8.22 2.12 ;
        RECT  8.00 1.84 8.16 3.48 ;
        RECT  7.10 1.84 7.26 3.48 ;
        RECT  6.90 1.84 7.26 2.12 ;
        RECT  6.06 1.84 6.22 3.48 ;
        RECT  5.86 1.84 6.22 2.12 ;
        RECT  0.38 2.48 0.66 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 11.60 0.28 ;
        RECT  11.08 -0.28 11.42 0.32 ;
        RECT  11.02 0.64 11.30 1.24 ;
        RECT  11.08 -0.28 11.24 1.24 ;
        RECT  9.98 0.64 10.26 1.24 ;
        RECT  10.04 -0.28 10.20 1.24 ;
        RECT  8.94 0.64 9.22 1.24 ;
        RECT  9.00 -0.28 9.16 1.24 ;
        RECT  7.94 0.88 8.22 1.16 ;
        RECT  8.00 -0.28 8.16 1.16 ;
        RECT  4.96 -0.28 5.24 0.72 ;
        RECT  0.38 -0.28 0.66 0.68 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  1.14 0.96 1.52 1.24 ;
        RECT  1.36 1.46 1.64 1.74 ;
        RECT  1.36 0.96 1.52 2.20 ;
        RECT  1.14 1.92 1.52 2.20 ;
        RECT  1.74 0.44 2.02 0.72 ;
        RECT  0.82 0.56 2.02 0.72 ;
        RECT  0.82 0.56 0.98 1.12 ;
        RECT  0.08 0.96 0.98 1.12 ;
        RECT  0.08 0.96 0.38 1.24 ;
        RECT  0.08 0.96 0.24 2.20 ;
        RECT  0.08 1.92 0.38 2.20 ;
        RECT  0.08 2.04 0.98 2.20 ;
        RECT  0.82 2.04 0.98 2.64 ;
        RECT  0.82 2.48 2.02 2.64 ;
        RECT  1.74 2.48 2.02 2.76 ;
        RECT  3.34 0.88 3.62 1.16 ;
        RECT  3.34 0.88 3.50 2.12 ;
        RECT  3.12 1.84 3.50 2.12 ;
        RECT  3.82 1.84 4.10 2.12 ;
        RECT  3.12 1.96 4.10 2.12 ;
        RECT  4.52 0.44 4.80 0.72 ;
        RECT  3.98 0.56 4.80 0.72 ;
        RECT  3.86 0.88 4.14 1.16 ;
        RECT  3.98 0.56 4.14 1.68 ;
        RECT  3.98 1.52 4.42 1.68 ;
        RECT  4.26 1.52 4.42 2.12 ;
        RECT  4.26 1.84 4.62 2.12 ;
        RECT  2.30 0.87 2.58 1.15 ;
        RECT  1.74 0.99 2.58 1.15 ;
        RECT  1.74 0.96 2.02 1.24 ;
        RECT  1.86 0.96 2.02 2.12 ;
        RECT  1.86 1.84 2.14 2.12 ;
        RECT  1.86 1.96 2.44 2.12 ;
        RECT  2.28 1.96 2.44 2.76 ;
        RECT  5.62 2.42 5.90 2.76 ;
        RECT  2.28 2.60 5.90 2.76 ;
        RECT  5.82 0.50 6.10 0.78 ;
        RECT  4.38 0.88 4.66 1.20 ;
        RECT  5.00 0.92 5.28 1.20 ;
        RECT  5.82 0.50 5.98 1.20 ;
        RECT  4.38 1.04 5.98 1.20 ;
        RECT  4.78 1.04 4.94 2.12 ;
        RECT  4.78 1.84 5.14 2.12 ;
        RECT  2.80 0.87 3.10 1.15 ;
        RECT  6.48 0.92 6.76 1.20 ;
        RECT  5.30 1.52 6.64 1.68 ;
        RECT  6.48 0.92 6.64 2.12 ;
        RECT  2.68 1.84 2.96 2.12 ;
        RECT  6.38 1.84 6.66 2.12 ;
        RECT  2.80 0.87 2.96 2.44 ;
        RECT  5.30 1.52 5.46 2.44 ;
        RECT  2.80 2.28 5.46 2.44 ;
        RECT  7.04 0.88 7.32 1.16 ;
        RECT  7.04 1.00 7.58 1.16 ;
        RECT  7.42 1.46 8.42 1.62 ;
        RECT  8.14 1.40 8.42 1.68 ;
        RECT  7.42 1.00 7.58 2.12 ;
        RECT  7.42 1.84 7.70 2.12 ;
        RECT  8.46 0.88 8.74 1.16 ;
        RECT  8.46 1.84 8.74 2.12 ;
        RECT  8.58 0.88 8.74 2.76 ;
        RECT  8.49 2.48 8.77 2.76 ;
    END
END DFFDRSP4V1_1

MACRO DFFDRSP4V1_0
    CLASS CORE ;
    FOREIGN DFFDRSP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 22.99  LAYER ME1  ;
        ANTENNADIFFAREA 10.06  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.21  LAYER ME1  ;
        ANTENNAMAXAREACAR 18.93  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.72 1.92 10.07 2.52 ;
        RECT  9.72 0.64 10.07 1.24 ;
        RECT  9.72 0.64 9.88 2.52 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 22.99  LAYER ME1  ;
        ANTENNADIFFAREA 10.18  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.21  LAYER ME1  ;
        ANTENNAMAXAREACAR 18.93  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.83 1.92 11.11 2.52 ;
        RECT  10.83 0.64 11.11 1.24 ;
        RECT  10.92 0.64 11.08 2.52 ;
        END
    END QB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.46 1.39 0.74 1.81 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.66 1.34 1.94 1.76 ;
        END
    END D
    PIN RB
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.42  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        ANTENNAMAXAREACAR 3.16  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.71 1.46 9.14 1.74 ;
        RECT  4.62 2.54 6.82 2.70 ;
        RECT  6.54 2.42 6.82 2.70 ;
        RECT  4.62 2.40 4.90 2.70 ;
        END
    END RB
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 12.00 3.48 ;
        RECT  11.41 2.88 11.82 3.48 ;
        RECT  11.35 1.92 11.63 2.52 ;
        RECT  11.41 1.92 11.57 3.48 ;
        RECT  10.31 1.92 10.59 2.52 ;
        RECT  10.38 1.92 10.54 3.48 ;
        RECT  9.27 1.92 9.55 2.52 ;
        RECT  9.33 1.92 9.49 3.48 ;
        RECT  8.77 1.90 9.05 2.18 ;
        RECT  8.83 1.90 8.99 3.48 ;
        RECT  7.73 1.90 8.01 2.18 ;
        RECT  7.79 1.90 7.95 3.48 ;
        RECT  3.76 2.08 5.08 2.24 ;
        RECT  4.80 1.96 5.08 2.24 ;
        RECT  4.30 2.08 4.46 3.48 ;
        RECT  3.76 1.96 4.04 2.24 ;
        RECT  1.64 1.92 1.92 2.20 ;
        RECT  1.72 1.92 1.88 3.48 ;
        RECT  0.62 1.97 0.90 2.25 ;
        RECT  0.68 1.97 0.84 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 12.00 0.28 ;
        RECT  11.41 -0.28 11.82 0.32 ;
        RECT  11.35 0.64 11.63 1.24 ;
        RECT  11.41 -0.28 11.57 1.24 ;
        RECT  10.31 0.64 10.59 1.24 ;
        RECT  10.37 -0.28 10.53 1.24 ;
        RECT  9.27 0.64 9.55 1.24 ;
        RECT  9.33 -0.28 9.49 1.24 ;
        RECT  7.75 0.96 8.03 1.24 ;
        RECT  7.82 -0.28 7.98 1.24 ;
        RECT  4.29 0.76 4.57 1.04 ;
        RECT  4.35 -0.28 4.51 1.04 ;
        RECT  1.64 0.76 1.92 1.04 ;
        RECT  1.70 -0.28 1.86 1.04 ;
        RECT  0.62 0.50 0.90 0.78 ;
        RECT  0.68 -0.28 0.84 0.78 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.07 0.50 0.38 0.78 ;
        RECT  0.07 0.94 1.16 1.10 ;
        RECT  0.88 0.94 1.16 1.22 ;
        RECT  0.07 0.50 0.23 2.25 ;
        RECT  0.07 1.97 0.38 2.25 ;
        RECT  1.14 0.50 1.48 0.78 ;
        RECT  1.14 1.97 1.48 2.25 ;
        RECT  1.32 0.50 1.48 2.70 ;
        RECT  1.28 2.42 1.56 2.70 ;
        RECT  2.16 0.76 2.44 1.04 ;
        RECT  2.22 0.76 2.38 2.20 ;
        RECT  2.16 1.92 2.44 2.20 ;
        RECT  3.20 0.76 3.48 1.04 ;
        RECT  3.26 0.76 3.42 2.20 ;
        RECT  3.20 1.92 3.48 2.20 ;
        RECT  3.32 1.92 3.48 2.62 ;
        RECT  3.32 2.46 4.00 2.62 ;
        RECT  3.72 2.46 4.00 2.74 ;
        RECT  2.80 0.44 3.94 0.60 ;
        RECT  2.80 0.44 2.96 1.04 ;
        RECT  2.68 0.76 2.96 1.04 ;
        RECT  3.78 0.44 3.94 1.36 ;
        RECT  3.78 1.20 5.08 1.36 ;
        RECT  4.80 1.20 5.08 1.48 ;
        RECT  2.74 0.76 2.90 2.20 ;
        RECT  2.68 1.92 2.96 2.20 ;
        RECT  5.04 0.76 5.40 1.04 ;
        RECT  3.59 1.52 3.87 1.80 ;
        RECT  3.59 1.64 5.40 1.80 ;
        RECT  5.24 0.76 5.40 2.24 ;
        RECT  5.24 1.96 5.60 2.24 ;
        RECT  5.76 0.44 7.37 0.60 ;
        RECT  7.09 0.44 7.37 0.72 ;
        RECT  5.56 0.76 5.92 1.04 ;
        RECT  5.76 0.44 5.92 2.24 ;
        RECT  5.76 1.96 6.12 2.24 ;
        RECT  6.69 1.90 6.97 2.24 ;
        RECT  5.76 2.08 6.97 2.24 ;
        RECT  6.08 0.76 6.36 1.12 ;
        RECT  6.08 0.96 7.51 1.12 ;
        RECT  7.21 0.96 7.51 1.24 ;
        RECT  6.21 0.96 6.37 1.81 ;
        RECT  6.21 1.53 6.49 1.81 ;
        RECT  7.21 0.96 7.37 2.18 ;
        RECT  7.21 1.90 7.49 2.18 ;
        RECT  8.79 0.44 9.07 0.72 ;
        RECT  8.33 0.96 8.95 1.12 ;
        RECT  8.79 0.44 8.95 1.24 ;
        RECT  8.65 0.96 8.95 1.24 ;
        RECT  7.55 1.52 8.49 1.68 ;
        RECT  7.55 1.46 7.83 1.74 ;
        RECT  8.33 0.96 8.49 2.18 ;
        RECT  8.25 1.90 8.53 2.18 ;
    END
END DFFDRSP4V1_0

MACRO DFFDRSP2V1_1
    CLASS CORE ;
    FOREIGN DFFDRSP2V1_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 20.58  LAYER ME1  ;
        ANTENNADIFFAREA 9.04  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.69  LAYER ME1  ;
        ANTENNAMAXAREACAR 29.78  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.06 1.46 10.32 1.74 ;
        RECT  9.98 1.90 10.26 2.50 ;
        RECT  10.06 0.64 10.26 2.50 ;
        RECT  9.98 0.64 10.26 1.24 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 20.58  LAYER ME1  ;
        ANTENNADIFFAREA 9.04  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.69  LAYER ME1  ;
        ANTENNAMAXAREACAR 29.78  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.06 1.46 9.54 1.74 ;
        RECT  8.94 1.90 9.22 2.50 ;
        RECT  9.06 0.64 9.22 2.50 ;
        RECT  8.94 0.64 9.22 1.24 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.40 0.72 1.76 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.88 1.40 1.20 1.76 ;
        END
    END CK
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.42 2.28 6.80 2.56 ;
        END
    END RB
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 10.40 0.28 ;
        RECT  9.94 -0.28 10.22 0.32 ;
        RECT  9.46 0.64 9.74 1.24 ;
        RECT  9.52 -0.28 9.68 1.24 ;
        RECT  7.94 0.88 8.22 1.16 ;
        RECT  8.00 -0.28 8.16 1.16 ;
        RECT  4.96 -0.28 5.24 0.72 ;
        RECT  0.38 -0.28 0.66 0.68 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 10.40 3.48 ;
        RECT  9.94 2.88 10.22 3.48 ;
        RECT  9.46 1.90 9.74 2.50 ;
        RECT  9.52 1.90 9.68 3.48 ;
        RECT  7.94 1.84 8.22 2.12 ;
        RECT  8.00 1.84 8.16 3.48 ;
        RECT  7.10 1.84 7.26 3.48 ;
        RECT  6.90 1.84 7.26 2.12 ;
        RECT  6.06 1.84 6.22 3.48 ;
        RECT  5.86 1.84 6.22 2.12 ;
        RECT  0.38 2.48 0.66 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  1.14 0.96 1.52 1.24 ;
        RECT  1.36 1.46 1.64 1.74 ;
        RECT  1.36 0.96 1.52 2.20 ;
        RECT  1.14 1.92 1.52 2.20 ;
        RECT  1.74 0.44 2.02 0.72 ;
        RECT  0.82 0.56 2.02 0.72 ;
        RECT  0.82 0.56 0.98 1.12 ;
        RECT  0.08 0.96 0.98 1.12 ;
        RECT  0.08 0.96 0.38 1.24 ;
        RECT  0.08 0.96 0.24 2.20 ;
        RECT  0.08 1.92 0.38 2.20 ;
        RECT  0.08 2.04 0.98 2.20 ;
        RECT  0.82 2.04 0.98 2.64 ;
        RECT  0.82 2.48 2.02 2.64 ;
        RECT  1.74 2.48 2.02 2.76 ;
        RECT  3.34 0.88 3.62 1.16 ;
        RECT  3.34 0.88 3.50 2.12 ;
        RECT  3.12 1.84 3.50 2.12 ;
        RECT  3.82 1.84 4.10 2.12 ;
        RECT  3.12 1.96 4.10 2.12 ;
        RECT  4.52 0.44 4.80 0.72 ;
        RECT  3.98 0.56 4.80 0.72 ;
        RECT  3.86 0.88 4.14 1.16 ;
        RECT  3.98 0.56 4.14 1.68 ;
        RECT  3.98 1.52 4.42 1.68 ;
        RECT  4.26 1.52 4.42 2.12 ;
        RECT  4.26 1.84 4.62 2.12 ;
        RECT  2.30 0.87 2.58 1.15 ;
        RECT  1.74 0.99 2.58 1.15 ;
        RECT  1.74 0.96 2.02 1.24 ;
        RECT  1.86 0.96 2.02 2.12 ;
        RECT  1.86 1.84 2.14 2.12 ;
        RECT  1.86 1.96 2.44 2.12 ;
        RECT  2.28 1.96 2.44 2.76 ;
        RECT  5.62 2.42 5.90 2.76 ;
        RECT  2.28 2.60 5.90 2.76 ;
        RECT  5.82 0.50 6.10 0.78 ;
        RECT  4.38 0.88 4.66 1.20 ;
        RECT  5.00 0.92 5.28 1.20 ;
        RECT  5.82 0.50 5.98 1.20 ;
        RECT  4.38 1.04 5.98 1.20 ;
        RECT  4.78 1.04 4.94 2.12 ;
        RECT  4.78 1.84 5.14 2.12 ;
        RECT  2.80 0.87 3.10 1.15 ;
        RECT  6.48 0.92 6.76 1.20 ;
        RECT  5.30 1.52 6.64 1.68 ;
        RECT  6.48 0.92 6.64 2.12 ;
        RECT  2.68 1.84 2.96 2.12 ;
        RECT  6.38 1.84 6.66 2.12 ;
        RECT  2.80 0.87 2.96 2.44 ;
        RECT  5.30 1.52 5.46 2.44 ;
        RECT  2.80 2.28 5.46 2.44 ;
        RECT  7.04 0.88 7.32 1.16 ;
        RECT  7.04 1.00 7.58 1.16 ;
        RECT  7.42 1.46 8.42 1.62 ;
        RECT  8.14 1.40 8.42 1.68 ;
        RECT  7.42 1.00 7.58 2.12 ;
        RECT  7.42 1.84 7.70 2.12 ;
        RECT  8.46 0.88 8.74 1.16 ;
        RECT  8.46 1.84 8.74 2.12 ;
        RECT  8.58 0.88 8.74 2.76 ;
        RECT  8.49 2.48 8.77 2.76 ;
    END
END DFFDRSP2V1_1

MACRO DFFDRSP2V1_0
    CLASS CORE ;
    FOREIGN DFFDRSP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN RB
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.42  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        ANTENNAMAXAREACAR 3.16  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.71 1.46 9.14 1.74 ;
        RECT  4.62 2.54 6.82 2.70 ;
        RECT  6.54 2.42 6.82 2.70 ;
        RECT  4.62 2.40 4.90 2.70 ;
        END
    END RB
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.66 1.34 1.94 1.76 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.46 1.39 0.74 1.81 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 20.76  LAYER ME1  ;
        ANTENNADIFFAREA 8.71  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.93  LAYER ME1  ;
        ANTENNAMAXAREACAR 22.41  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.31 1.92 10.68 2.52 ;
        RECT  10.52 0.64 10.68 2.52 ;
        RECT  10.31 0.64 10.68 1.24 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 20.76  LAYER ME1  ;
        ANTENNADIFFAREA 8.71  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.93  LAYER ME1  ;
        ANTENNAMAXAREACAR 22.41  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.27 1.92 9.55 2.52 ;
        RECT  9.27 0.64 9.55 1.24 ;
        RECT  9.32 0.64 9.48 2.52 ;
        END
    END Q
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 10.80 0.28 ;
        RECT  10.34 -0.28 10.62 0.32 ;
        RECT  9.79 0.64 10.07 1.24 ;
        RECT  9.85 -0.28 10.01 1.24 ;
        RECT  7.75 0.96 8.03 1.24 ;
        RECT  7.82 -0.28 7.98 1.24 ;
        RECT  4.29 0.76 4.57 1.04 ;
        RECT  4.35 -0.28 4.51 1.04 ;
        RECT  1.64 0.76 1.92 1.04 ;
        RECT  1.70 -0.28 1.86 1.04 ;
        RECT  0.62 0.50 0.90 0.78 ;
        RECT  0.68 -0.28 0.84 0.78 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 10.80 3.48 ;
        RECT  10.34 2.88 10.62 3.48 ;
        RECT  9.79 1.92 10.07 2.52 ;
        RECT  9.85 1.92 10.01 3.48 ;
        RECT  8.77 1.90 9.05 2.18 ;
        RECT  8.83 1.90 8.99 3.48 ;
        RECT  7.73 1.90 8.01 2.18 ;
        RECT  7.79 1.90 7.95 3.48 ;
        RECT  3.76 2.08 5.08 2.24 ;
        RECT  4.80 1.96 5.08 2.24 ;
        RECT  4.30 2.08 4.46 3.48 ;
        RECT  3.76 1.96 4.04 2.24 ;
        RECT  1.64 1.92 1.92 2.20 ;
        RECT  1.72 1.92 1.88 3.48 ;
        RECT  0.62 1.97 0.90 2.25 ;
        RECT  0.68 1.97 0.84 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.07 0.50 0.38 0.78 ;
        RECT  0.07 0.94 1.16 1.10 ;
        RECT  0.88 0.94 1.16 1.22 ;
        RECT  0.07 0.50 0.23 2.25 ;
        RECT  0.07 1.97 0.38 2.25 ;
        RECT  1.14 0.50 1.48 0.78 ;
        RECT  1.14 1.97 1.48 2.25 ;
        RECT  1.32 0.50 1.48 2.70 ;
        RECT  1.28 2.42 1.56 2.70 ;
        RECT  2.16 0.76 2.44 1.04 ;
        RECT  2.22 0.76 2.38 2.20 ;
        RECT  2.16 1.92 2.44 2.20 ;
        RECT  3.20 0.76 3.48 1.04 ;
        RECT  3.26 0.76 3.42 2.20 ;
        RECT  3.20 1.92 3.48 2.20 ;
        RECT  3.32 1.92 3.48 2.62 ;
        RECT  3.32 2.46 4.00 2.62 ;
        RECT  3.72 2.46 4.00 2.74 ;
        RECT  2.80 0.44 3.94 0.60 ;
        RECT  2.80 0.44 2.96 1.04 ;
        RECT  2.68 0.76 2.96 1.04 ;
        RECT  3.78 0.44 3.94 1.36 ;
        RECT  3.78 1.20 5.08 1.36 ;
        RECT  4.80 1.20 5.08 1.48 ;
        RECT  2.74 0.76 2.90 2.20 ;
        RECT  2.68 1.92 2.96 2.20 ;
        RECT  5.04 0.76 5.40 1.04 ;
        RECT  3.59 1.52 3.87 1.80 ;
        RECT  3.59 1.64 5.40 1.80 ;
        RECT  5.24 0.76 5.40 2.24 ;
        RECT  5.24 1.96 5.60 2.24 ;
        RECT  5.76 0.44 7.37 0.60 ;
        RECT  7.09 0.44 7.37 0.72 ;
        RECT  5.56 0.76 5.92 1.04 ;
        RECT  5.76 0.44 5.92 2.24 ;
        RECT  5.76 1.96 6.12 2.24 ;
        RECT  6.69 1.90 6.97 2.24 ;
        RECT  5.76 2.08 6.97 2.24 ;
        RECT  6.08 0.76 6.36 1.12 ;
        RECT  6.08 0.96 7.51 1.12 ;
        RECT  7.21 0.96 7.51 1.24 ;
        RECT  6.21 0.96 6.37 1.81 ;
        RECT  6.21 1.53 6.49 1.81 ;
        RECT  7.21 0.96 7.37 2.18 ;
        RECT  7.21 1.90 7.49 2.18 ;
        RECT  8.79 0.44 9.07 0.72 ;
        RECT  8.33 0.96 8.95 1.12 ;
        RECT  8.79 0.44 8.95 1.24 ;
        RECT  8.65 0.96 8.95 1.24 ;
        RECT  7.55 1.52 8.49 1.68 ;
        RECT  7.55 1.46 7.83 1.74 ;
        RECT  8.33 0.96 8.49 2.18 ;
        RECT  8.25 1.90 8.53 2.18 ;
    END
END DFFDRSP2V1_0

MACRO DFFDRSP1V1_1
    CLASS CORE ;
    FOREIGN DFFDRSP1V1_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.40 0.72 1.76 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.88 1.40 1.20 1.76 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 19.84  LAYER ME1  ;
        ANTENNADIFFAREA 8.34  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.54  LAYER ME1  ;
        ANTENNAMAXAREACAR 36.91  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.06 1.46 10.32 1.74 ;
        RECT  9.98 1.90 10.26 2.18 ;
        RECT  10.06 0.88 10.26 2.18 ;
        RECT  9.98 0.88 10.26 1.16 ;
        END
    END QB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.42 2.28 6.80 2.56 ;
        END
    END RB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 20.16  LAYER ME1  ;
        ANTENNADIFFAREA 8.34  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.54  LAYER ME1  ;
        ANTENNAMAXAREACAR 37.50  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.06 1.46 9.54 1.74 ;
        RECT  8.94 1.90 9.22 2.18 ;
        RECT  9.06 0.88 9.22 2.18 ;
        RECT  8.94 0.88 9.22 1.16 ;
        END
    END Q
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 10.40 3.48 ;
        RECT  9.94 2.88 10.22 3.48 ;
        RECT  9.46 1.90 9.74 2.18 ;
        RECT  9.52 1.90 9.68 3.48 ;
        RECT  7.94 1.84 8.22 2.12 ;
        RECT  8.00 1.84 8.16 3.48 ;
        RECT  7.10 1.84 7.26 3.48 ;
        RECT  6.90 1.84 7.26 2.12 ;
        RECT  6.06 1.84 6.22 3.48 ;
        RECT  5.86 1.84 6.22 2.12 ;
        RECT  0.38 2.48 0.66 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 10.40 0.28 ;
        RECT  9.94 -0.28 10.22 0.32 ;
        RECT  9.46 0.88 9.74 1.16 ;
        RECT  9.52 -0.28 9.68 1.16 ;
        RECT  7.94 0.88 8.22 1.16 ;
        RECT  8.00 -0.28 8.16 1.16 ;
        RECT  4.96 -0.28 5.24 0.72 ;
        RECT  0.38 -0.28 0.66 0.68 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  1.14 0.96 1.52 1.24 ;
        RECT  1.36 1.46 1.64 1.74 ;
        RECT  1.36 0.96 1.52 2.20 ;
        RECT  1.14 1.92 1.52 2.20 ;
        RECT  1.74 0.44 2.02 0.72 ;
        RECT  0.82 0.56 2.02 0.72 ;
        RECT  0.82 0.56 0.98 1.12 ;
        RECT  0.08 0.96 0.98 1.12 ;
        RECT  0.08 0.96 0.38 1.24 ;
        RECT  0.08 0.96 0.24 2.20 ;
        RECT  0.08 1.92 0.38 2.20 ;
        RECT  0.08 2.04 0.98 2.20 ;
        RECT  0.82 2.04 0.98 2.64 ;
        RECT  0.82 2.48 2.02 2.64 ;
        RECT  1.74 2.48 2.02 2.76 ;
        RECT  3.34 0.88 3.62 1.16 ;
        RECT  3.34 0.88 3.50 2.12 ;
        RECT  3.12 1.84 3.50 2.12 ;
        RECT  3.82 1.84 4.10 2.12 ;
        RECT  3.12 1.96 4.10 2.12 ;
        RECT  4.52 0.44 4.80 0.72 ;
        RECT  3.98 0.56 4.80 0.72 ;
        RECT  3.86 0.88 4.14 1.16 ;
        RECT  3.98 0.56 4.14 1.68 ;
        RECT  3.98 1.52 4.42 1.68 ;
        RECT  4.26 1.52 4.42 2.12 ;
        RECT  4.26 1.84 4.62 2.12 ;
        RECT  2.30 0.87 2.58 1.15 ;
        RECT  1.74 0.99 2.58 1.15 ;
        RECT  1.74 0.96 2.02 1.24 ;
        RECT  1.86 0.96 2.02 2.12 ;
        RECT  1.86 1.84 2.14 2.12 ;
        RECT  1.86 1.96 2.44 2.12 ;
        RECT  2.28 1.96 2.44 2.76 ;
        RECT  5.62 2.42 5.90 2.76 ;
        RECT  2.28 2.60 5.90 2.76 ;
        RECT  5.82 0.50 6.10 0.78 ;
        RECT  4.38 0.88 4.66 1.20 ;
        RECT  5.00 0.92 5.28 1.20 ;
        RECT  5.82 0.50 5.98 1.20 ;
        RECT  4.38 1.04 5.98 1.20 ;
        RECT  4.78 1.04 4.94 2.12 ;
        RECT  4.78 1.84 5.14 2.12 ;
        RECT  2.80 0.87 3.10 1.15 ;
        RECT  6.48 0.92 6.76 1.20 ;
        RECT  5.30 1.52 6.64 1.68 ;
        RECT  6.48 0.92 6.64 2.12 ;
        RECT  2.68 1.84 2.96 2.12 ;
        RECT  6.38 1.84 6.66 2.12 ;
        RECT  2.80 0.87 2.96 2.44 ;
        RECT  5.30 1.52 5.46 2.44 ;
        RECT  2.80 2.28 5.46 2.44 ;
        RECT  7.04 0.88 7.32 1.16 ;
        RECT  7.04 1.00 7.58 1.16 ;
        RECT  7.42 1.46 8.42 1.62 ;
        RECT  8.14 1.40 8.42 1.68 ;
        RECT  7.42 1.00 7.58 2.12 ;
        RECT  7.42 1.84 7.70 2.12 ;
        RECT  8.46 0.88 8.74 1.16 ;
        RECT  8.46 1.84 8.74 2.12 ;
        RECT  8.58 0.88 8.74 2.76 ;
        RECT  8.49 2.48 8.77 2.76 ;
    END
END DFFDRSP1V1_1

MACRO DFFDRSP1V1_0
    CLASS CORE ;
    FOREIGN DFFDRSP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 19.14  LAYER ME1  ;
        ANTENNADIFFAREA 7.84  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.54  LAYER ME1  ;
        ANTENNAMAXAREACAR 35.61  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.77 1.92 10.05 2.20 ;
        RECT  9.77 0.75 10.05 1.03 ;
        RECT  9.77 0.75 9.93 2.20 ;
        RECT  9.66 1.46 9.93 1.74 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 19.47  LAYER ME1  ;
        ANTENNADIFFAREA 7.84  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.54  LAYER ME1  ;
        ANTENNAMAXAREACAR 36.22  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.85 1.46 9.14 1.74 ;
        RECT  8.73 1.92 9.01 2.20 ;
        RECT  8.85 0.75 9.01 2.20 ;
        RECT  8.73 0.75 9.01 1.03 ;
        END
    END QB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.88 1.34 1.16 1.76 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.34 0.72 1.76 ;
        END
    END D
    PIN RB
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.42  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        ANTENNAMAXAREACAR 3.16  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.06 1.46 8.49 1.74 ;
        RECT  4.08 2.54 6.28 2.70 ;
        RECT  6.00 2.42 6.28 2.70 ;
        RECT  4.08 2.40 4.36 2.70 ;
        END
    END RB
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 10.40 0.28 ;
        RECT  9.94 -0.28 10.22 0.32 ;
        RECT  9.25 0.75 9.53 1.03 ;
        RECT  9.31 -0.28 9.47 1.03 ;
        RECT  7.21 0.96 7.49 1.24 ;
        RECT  7.28 -0.28 7.44 1.24 ;
        RECT  3.77 0.76 4.05 1.04 ;
        RECT  3.83 -0.28 3.99 1.04 ;
        RECT  0.62 0.76 0.90 1.04 ;
        RECT  0.69 -0.28 0.85 1.04 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 10.40 3.48 ;
        RECT  9.94 2.88 10.22 3.48 ;
        RECT  9.25 1.92 9.53 2.20 ;
        RECT  9.31 1.92 9.47 3.48 ;
        RECT  8.23 1.90 8.51 2.18 ;
        RECT  8.29 1.90 8.45 3.48 ;
        RECT  7.19 1.90 7.47 2.18 ;
        RECT  7.25 1.90 7.41 3.48 ;
        RECT  3.22 2.08 4.54 2.24 ;
        RECT  4.26 1.96 4.54 2.24 ;
        RECT  3.76 2.08 3.92 3.48 ;
        RECT  3.22 1.96 3.50 2.24 ;
        RECT  0.38 2.48 0.66 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  1.14 0.76 1.48 1.04 ;
        RECT  1.32 1.21 1.64 1.49 ;
        RECT  1.32 0.76 1.48 2.20 ;
        RECT  1.14 1.92 1.48 2.20 ;
        RECT  0.08 0.76 0.38 1.04 ;
        RECT  1.64 0.76 1.96 1.04 ;
        RECT  0.08 0.76 0.24 2.20 ;
        RECT  0.08 1.92 0.38 2.20 ;
        RECT  0.08 2.04 0.98 2.20 ;
        RECT  1.80 0.76 1.96 2.20 ;
        RECT  0.82 2.04 0.98 2.52 ;
        RECT  1.64 1.92 1.80 2.52 ;
        RECT  0.82 2.36 1.80 2.52 ;
        RECT  2.68 0.76 2.96 1.04 ;
        RECT  2.72 0.76 2.88 2.20 ;
        RECT  2.68 1.92 2.96 2.20 ;
        RECT  2.80 1.92 2.96 2.62 ;
        RECT  2.80 2.46 3.46 2.62 ;
        RECT  3.18 2.46 3.46 2.74 ;
        RECT  2.26 0.44 3.40 0.60 ;
        RECT  2.26 0.44 2.42 1.04 ;
        RECT  2.16 0.76 2.44 1.04 ;
        RECT  3.24 0.44 3.40 1.36 ;
        RECT  3.24 1.20 4.54 1.36 ;
        RECT  4.26 1.20 4.54 1.48 ;
        RECT  2.20 0.76 2.36 2.20 ;
        RECT  2.16 1.92 2.44 2.20 ;
        RECT  4.50 0.76 4.86 1.04 ;
        RECT  3.07 1.52 3.35 1.80 ;
        RECT  3.07 1.64 4.86 1.80 ;
        RECT  4.70 0.76 4.86 2.24 ;
        RECT  4.70 1.96 5.06 2.24 ;
        RECT  5.22 0.44 6.83 0.60 ;
        RECT  6.55 0.44 6.83 0.72 ;
        RECT  5.02 0.76 5.38 1.04 ;
        RECT  5.22 0.44 5.38 2.24 ;
        RECT  5.22 1.96 5.58 2.24 ;
        RECT  6.15 1.90 6.43 2.24 ;
        RECT  5.22 2.08 6.43 2.24 ;
        RECT  5.54 0.76 5.82 1.12 ;
        RECT  5.54 0.96 6.97 1.12 ;
        RECT  6.67 0.96 6.97 1.24 ;
        RECT  5.67 0.96 5.83 1.81 ;
        RECT  5.67 1.53 5.95 1.81 ;
        RECT  6.67 0.96 6.83 2.18 ;
        RECT  6.67 1.90 6.95 2.18 ;
        RECT  8.25 0.44 8.53 0.72 ;
        RECT  7.74 0.96 8.41 1.12 ;
        RECT  8.25 0.44 8.41 1.24 ;
        RECT  8.11 0.96 8.41 1.24 ;
        RECT  7.01 1.52 7.90 1.68 ;
        RECT  7.01 1.46 7.29 1.74 ;
        RECT  7.74 0.96 7.90 2.18 ;
        RECT  7.71 1.90 7.99 2.18 ;
    END
END DFFDRSP1V1_0

MACRO DFFDRHZSP8V1_0
    CLASS CORE ;
    FOREIGN DFFDRHZSP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 17.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.43  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  16.77 1.46 17.17 1.74 ;
        END
    END E
    PIN QZ
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 33.31  LAYER ME1  ;
        ANTENNADIFFAREA 16.14  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.48  LAYER ME1  ;
        ANTENNAMAXAREACAR 22.53  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  15.43 1.90 15.71 2.18 ;
        RECT  15.43 0.96 15.71 1.24 ;
        RECT  15.43 0.96 15.59 2.18 ;
        RECT  14.46 1.52 15.59 1.68 ;
        RECT  14.46 1.46 14.75 1.74 ;
        RECT  14.39 1.90 14.67 2.18 ;
        RECT  14.46 0.96 14.67 2.18 ;
        RECT  14.39 0.96 14.67 1.24 ;
        END
    END QZ
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 33.31  LAYER ME1  ;
        ANTENNADIFFAREA 16.37  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.48  LAYER ME1  ;
        ANTENNAMAXAREACAR 22.53  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.83 1.90 13.11 2.50 ;
        RECT  12.83 0.64 13.11 1.24 ;
        RECT  12.83 0.64 12.99 2.50 ;
        RECT  11.66 1.52 12.99 1.68 ;
        RECT  11.79 1.90 12.07 2.50 ;
        RECT  11.79 0.64 12.07 1.24 ;
        RECT  11.79 0.64 11.95 2.50 ;
        RECT  11.66 1.46 11.95 1.74 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.20  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.83  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.81 1.19 2.25 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  0.91 0.81 1.19 1.09 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.22 1.40 3.54 1.76 ;
        END
    END CK
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.79 2.28 9.17 2.56 ;
        END
    END RB
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.87  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 12.90  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.06 1.46 2.34 1.74 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.81 2.23 2.25 ;
        RECT  1.95 0.81 2.23 1.09 ;
        END
    END TD
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END SEL
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 17.60 0.28 ;
        RECT  17.01 -0.28 17.42 0.32 ;
        RECT  16.95 0.64 17.23 1.24 ;
        RECT  17.01 -0.28 17.17 1.24 ;
        RECT  13.35 0.64 13.63 1.24 ;
        RECT  13.41 -0.28 13.57 1.24 ;
        RECT  12.31 0.64 12.59 1.24 ;
        RECT  12.37 -0.28 12.53 1.24 ;
        RECT  11.27 0.64 11.55 1.24 ;
        RECT  11.33 -0.28 11.49 1.24 ;
        RECT  10.27 0.88 10.55 1.16 ;
        RECT  10.33 -0.28 10.49 1.16 ;
        RECT  7.29 -0.28 7.57 0.72 ;
        RECT  2.71 -0.28 2.99 0.68 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 17.60 3.48 ;
        RECT  17.01 2.88 17.42 3.48 ;
        RECT  16.95 1.90 17.23 2.50 ;
        RECT  17.01 1.90 17.17 3.48 ;
        RECT  13.35 1.90 13.63 2.50 ;
        RECT  13.41 1.90 13.57 3.48 ;
        RECT  12.31 1.90 12.59 2.50 ;
        RECT  12.37 1.90 12.53 3.48 ;
        RECT  11.27 1.90 11.55 2.50 ;
        RECT  11.33 1.90 11.49 3.48 ;
        RECT  10.27 1.84 10.55 2.12 ;
        RECT  10.33 1.84 10.49 3.48 ;
        RECT  9.43 1.84 9.59 3.48 ;
        RECT  9.23 1.84 9.59 2.12 ;
        RECT  8.39 1.84 8.55 3.48 ;
        RECT  8.19 1.84 8.55 2.12 ;
        RECT  2.71 2.52 2.99 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  1.55 1.97 1.71 2.57 ;
        RECT  1.55 2.41 2.37 2.57 ;
        RECT  2.09 2.41 2.37 2.69 ;
        RECT  3.47 0.96 3.86 1.24 ;
        RECT  3.70 1.46 4.02 1.74 ;
        RECT  3.70 0.96 3.86 2.20 ;
        RECT  3.47 1.92 3.86 2.20 ;
        RECT  4.07 0.44 4.35 0.72 ;
        RECT  3.15 0.56 4.35 0.72 ;
        RECT  3.15 0.56 3.31 1.12 ;
        RECT  2.43 0.96 3.31 1.12 ;
        RECT  2.43 0.96 2.71 1.24 ;
        RECT  2.55 0.96 2.71 2.20 ;
        RECT  2.43 1.92 2.71 2.20 ;
        RECT  2.43 2.04 3.31 2.20 ;
        RECT  3.15 2.04 3.31 2.64 ;
        RECT  3.15 2.48 4.35 2.64 ;
        RECT  4.07 2.48 4.35 2.76 ;
        RECT  5.67 0.88 5.95 1.16 ;
        RECT  5.67 0.88 5.83 2.12 ;
        RECT  5.45 1.84 5.83 2.12 ;
        RECT  6.15 1.84 6.43 2.12 ;
        RECT  5.45 1.96 6.43 2.12 ;
        RECT  6.85 0.44 7.13 0.72 ;
        RECT  6.31 0.56 7.13 0.72 ;
        RECT  6.19 0.88 6.47 1.16 ;
        RECT  6.31 0.56 6.47 1.68 ;
        RECT  6.31 1.52 6.75 1.68 ;
        RECT  6.59 1.52 6.75 2.12 ;
        RECT  6.59 1.84 6.95 2.12 ;
        RECT  4.63 0.87 4.91 1.15 ;
        RECT  4.07 0.99 4.91 1.15 ;
        RECT  4.07 0.96 4.35 1.24 ;
        RECT  4.19 0.96 4.35 2.12 ;
        RECT  4.19 1.84 4.47 2.12 ;
        RECT  4.19 1.96 4.77 2.12 ;
        RECT  4.61 1.96 4.77 2.76 ;
        RECT  7.95 2.42 8.23 2.76 ;
        RECT  4.61 2.60 8.23 2.76 ;
        RECT  8.15 0.50 8.43 0.78 ;
        RECT  6.71 0.88 6.99 1.20 ;
        RECT  7.33 0.92 7.61 1.20 ;
        RECT  8.15 0.50 8.31 1.20 ;
        RECT  6.71 1.04 8.31 1.20 ;
        RECT  7.11 1.04 7.27 2.12 ;
        RECT  7.11 1.84 7.47 2.12 ;
        RECT  5.13 0.87 5.43 1.15 ;
        RECT  8.81 0.92 9.09 1.20 ;
        RECT  7.63 1.52 8.97 1.68 ;
        RECT  8.81 0.92 8.97 2.12 ;
        RECT  5.01 1.84 5.29 2.12 ;
        RECT  8.71 1.84 8.99 2.12 ;
        RECT  5.13 0.87 5.29 2.44 ;
        RECT  7.63 1.52 7.79 2.44 ;
        RECT  5.13 2.28 7.79 2.44 ;
        RECT  9.37 0.88 9.65 1.16 ;
        RECT  9.37 1.00 9.91 1.16 ;
        RECT  9.75 1.46 10.75 1.62 ;
        RECT  10.47 1.40 10.75 1.68 ;
        RECT  9.75 1.00 9.91 2.12 ;
        RECT  9.75 1.84 10.03 2.12 ;
        RECT  10.79 0.88 11.07 1.16 ;
        RECT  10.79 1.84 11.07 2.12 ;
        RECT  10.91 0.88 11.07 2.76 ;
        RECT  10.82 2.48 11.10 2.76 ;
        RECT  13.87 1.90 14.15 2.50 ;
        RECT  14.91 1.90 15.19 2.50 ;
        RECT  15.95 1.90 16.23 2.50 ;
        RECT  13.87 2.34 16.23 2.50 ;
        RECT  13.87 0.64 16.23 0.80 ;
        RECT  13.87 0.64 14.15 1.24 ;
        RECT  14.91 0.64 15.19 1.24 ;
        RECT  15.95 0.64 16.23 1.24 ;
        RECT  16.43 0.64 16.71 1.24 ;
        RECT  16.29 1.46 16.59 1.74 ;
        RECT  16.43 0.64 16.59 2.50 ;
        RECT  16.43 1.90 16.71 2.50 ;
    END
END DFFDRHZSP8V1_0

MACRO DFFDRHZSP4V1_0
    CLASS CORE ;
    FOREIGN DFFDRHZSP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.22 1.40 3.54 1.76 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 28.99  LAYER ME1  ;
        ANTENNADIFFAREA 13.43  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.05  LAYER ME1  ;
        ANTENNAMAXAREACAR 27.71  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.79 1.90 12.07 2.50 ;
        RECT  11.79 0.64 12.07 1.24 ;
        RECT  11.79 0.64 11.95 2.50 ;
        RECT  11.66 1.46 11.95 1.74 ;
        END
    END Q
    PIN QZ
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 28.69  LAYER ME1  ;
        ANTENNADIFFAREA 13.45  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.05  LAYER ME1  ;
        ANTENNAMAXAREACAR 27.41  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.35 1.90 13.63 2.18 ;
        RECT  13.35 0.96 13.63 1.24 ;
        RECT  13.35 0.96 13.54 2.18 ;
        RECT  13.26 1.46 13.54 1.74 ;
        END
    END QZ
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.26  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.69 1.46 15.14 1.74 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.20  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.83  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.81 1.19 2.25 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  0.91 0.81 1.19 1.09 ;
        END
    END D
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END SEL
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.87  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 12.90  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.06 1.46 2.34 1.74 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.81 2.23 2.25 ;
        RECT  1.95 0.81 2.23 1.09 ;
        END
    END TD
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.79 2.28 9.17 2.56 ;
        END
    END RB
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 15.60 0.28 ;
        RECT  14.98 -0.28 15.42 0.32 ;
        RECT  14.87 0.74 15.15 1.24 ;
        RECT  14.98 -0.28 15.14 1.24 ;
        RECT  12.31 0.64 12.59 1.24 ;
        RECT  12.37 -0.28 12.53 1.24 ;
        RECT  11.27 0.64 11.55 1.24 ;
        RECT  11.33 -0.28 11.49 1.24 ;
        RECT  10.27 0.88 10.55 1.16 ;
        RECT  10.33 -0.28 10.49 1.16 ;
        RECT  7.29 -0.28 7.57 0.72 ;
        RECT  2.71 -0.28 2.99 0.68 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 15.60 3.48 ;
        RECT  14.98 2.88 15.42 3.48 ;
        RECT  14.87 1.90 15.15 2.40 ;
        RECT  14.98 1.90 15.14 3.48 ;
        RECT  12.31 1.90 12.59 2.50 ;
        RECT  12.37 1.90 12.53 3.48 ;
        RECT  11.27 1.90 11.55 2.50 ;
        RECT  11.33 1.90 11.49 3.48 ;
        RECT  10.27 1.84 10.55 2.12 ;
        RECT  10.33 1.84 10.49 3.48 ;
        RECT  9.43 1.84 9.59 3.48 ;
        RECT  9.23 1.84 9.59 2.12 ;
        RECT  8.39 1.84 8.55 3.48 ;
        RECT  8.19 1.84 8.55 2.12 ;
        RECT  2.71 2.52 2.99 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  1.55 1.97 1.71 2.57 ;
        RECT  1.55 2.41 2.37 2.57 ;
        RECT  2.09 2.41 2.37 2.69 ;
        RECT  3.47 0.96 3.86 1.24 ;
        RECT  3.70 1.46 4.02 1.74 ;
        RECT  3.70 0.96 3.86 2.20 ;
        RECT  3.47 1.92 3.86 2.20 ;
        RECT  4.07 0.44 4.35 0.72 ;
        RECT  3.15 0.56 4.35 0.72 ;
        RECT  3.15 0.56 3.31 1.12 ;
        RECT  2.43 0.96 3.31 1.12 ;
        RECT  2.43 0.96 2.71 1.24 ;
        RECT  2.55 0.96 2.71 2.20 ;
        RECT  2.43 1.92 2.71 2.20 ;
        RECT  2.43 2.04 3.31 2.20 ;
        RECT  3.15 2.04 3.31 2.64 ;
        RECT  3.15 2.48 4.35 2.64 ;
        RECT  4.07 2.48 4.35 2.76 ;
        RECT  5.67 0.88 5.95 1.16 ;
        RECT  5.67 0.88 5.83 2.12 ;
        RECT  5.45 1.84 5.83 2.12 ;
        RECT  6.15 1.84 6.43 2.12 ;
        RECT  5.45 1.96 6.43 2.12 ;
        RECT  6.85 0.44 7.13 0.72 ;
        RECT  6.31 0.56 7.13 0.72 ;
        RECT  6.19 0.88 6.47 1.16 ;
        RECT  6.31 0.56 6.47 1.68 ;
        RECT  6.31 1.52 6.75 1.68 ;
        RECT  6.59 1.52 6.75 2.12 ;
        RECT  6.59 1.84 6.95 2.12 ;
        RECT  4.63 0.87 4.91 1.15 ;
        RECT  4.07 0.99 4.91 1.15 ;
        RECT  4.07 0.96 4.35 1.24 ;
        RECT  4.19 0.96 4.35 2.12 ;
        RECT  4.19 1.84 4.47 2.12 ;
        RECT  4.19 1.96 4.77 2.12 ;
        RECT  4.61 1.96 4.77 2.76 ;
        RECT  7.95 2.42 8.23 2.76 ;
        RECT  4.61 2.60 8.23 2.76 ;
        RECT  8.15 0.50 8.43 0.78 ;
        RECT  6.71 0.88 6.99 1.20 ;
        RECT  7.33 0.92 7.61 1.20 ;
        RECT  8.15 0.50 8.31 1.20 ;
        RECT  6.71 1.04 8.31 1.20 ;
        RECT  7.11 1.04 7.27 2.12 ;
        RECT  7.11 1.84 7.47 2.12 ;
        RECT  5.13 0.87 5.43 1.15 ;
        RECT  8.81 0.92 9.09 1.20 ;
        RECT  7.63 1.52 8.97 1.68 ;
        RECT  8.81 0.92 8.97 2.12 ;
        RECT  5.01 1.84 5.29 2.12 ;
        RECT  8.71 1.84 8.99 2.12 ;
        RECT  5.13 0.87 5.29 2.44 ;
        RECT  7.63 1.52 7.79 2.44 ;
        RECT  5.13 2.28 7.79 2.44 ;
        RECT  9.37 0.88 9.65 1.16 ;
        RECT  9.37 1.00 9.91 1.16 ;
        RECT  9.75 1.46 10.75 1.62 ;
        RECT  10.47 1.40 10.75 1.68 ;
        RECT  9.75 1.00 9.91 2.12 ;
        RECT  9.75 1.84 10.03 2.12 ;
        RECT  10.79 0.88 11.07 1.16 ;
        RECT  10.79 1.84 11.07 2.12 ;
        RECT  10.91 0.88 11.07 2.76 ;
        RECT  10.82 2.48 11.10 2.76 ;
        RECT  12.83 1.90 13.11 2.50 ;
        RECT  13.87 1.90 14.15 2.50 ;
        RECT  12.83 2.34 14.15 2.50 ;
        RECT  12.83 0.64 14.15 0.80 ;
        RECT  12.83 0.64 13.11 1.24 ;
        RECT  13.87 0.64 14.15 1.24 ;
        RECT  14.35 0.74 14.63 1.24 ;
        RECT  14.21 1.46 14.51 1.74 ;
        RECT  14.35 0.74 14.51 2.40 ;
        RECT  14.35 1.90 14.63 2.40 ;
    END
END DFFDRHZSP4V1_0

MACRO DFFDRHZSP2V1_0
    CLASS CORE ;
    FOREIGN DFFDRHZSP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.17  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.49 1.46 13.94 1.74 ;
        END
    END E
    PIN QZ
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 26.43  LAYER ME1  ;
        ANTENNADIFFAREA 11.54  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.83  LAYER ME1  ;
        ANTENNAMAXAREACAR 31.83  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.69 1.90 12.97 2.50 ;
        RECT  12.69 0.64 12.97 1.24 ;
        RECT  12.69 0.64 12.85 2.50 ;
        RECT  12.46 1.46 12.85 1.74 ;
        END
    END QZ
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 26.43  LAYER ME1  ;
        ANTENNADIFFAREA 11.54  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.83  LAYER ME1  ;
        ANTENNAMAXAREACAR 31.83  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.27 1.90 11.55 2.50 ;
        RECT  11.27 0.64 11.55 1.24 ;
        RECT  11.27 0.64 11.54 2.50 ;
        RECT  11.26 1.46 11.54 1.74 ;
        END
    END Q
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.75 2.28 9.13 2.56 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.22 1.40 3.54 1.76 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.87  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 12.90  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.06 1.46 2.34 1.74 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.81 2.23 2.25 ;
        RECT  1.95 0.81 2.23 1.09 ;
        END
    END TD
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END SEL
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.20  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.83  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.81 1.19 2.25 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  0.91 0.81 1.19 1.09 ;
        END
    END D
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 14.40 0.28 ;
        RECT  13.78 -0.28 14.22 0.32 ;
        RECT  13.69 0.84 13.97 1.24 ;
        RECT  13.78 -0.28 13.94 1.24 ;
        RECT  11.79 0.64 12.07 1.24 ;
        RECT  11.85 -0.28 12.01 1.24 ;
        RECT  10.27 0.88 10.55 1.16 ;
        RECT  10.33 -0.28 10.49 1.16 ;
        RECT  7.29 -0.28 7.57 0.72 ;
        RECT  2.71 -0.28 2.99 0.68 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 14.40 3.48 ;
        RECT  13.78 2.88 14.22 3.48 ;
        RECT  13.69 1.90 13.97 2.30 ;
        RECT  13.78 1.90 13.94 3.48 ;
        RECT  11.79 1.90 12.07 2.50 ;
        RECT  11.85 1.90 12.01 3.48 ;
        RECT  10.27 1.84 10.55 2.12 ;
        RECT  10.33 1.84 10.49 3.48 ;
        RECT  9.43 1.84 9.59 3.48 ;
        RECT  9.23 1.84 9.59 2.12 ;
        RECT  8.39 1.84 8.55 3.48 ;
        RECT  8.19 1.84 8.55 2.12 ;
        RECT  2.71 2.52 2.99 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  1.55 1.97 1.71 2.57 ;
        RECT  1.55 2.41 2.37 2.57 ;
        RECT  2.09 2.41 2.37 2.69 ;
        RECT  3.47 0.96 3.86 1.24 ;
        RECT  3.70 1.46 4.02 1.74 ;
        RECT  3.70 0.96 3.86 2.20 ;
        RECT  3.47 1.92 3.86 2.20 ;
        RECT  4.07 0.44 4.35 0.72 ;
        RECT  3.15 0.56 4.35 0.72 ;
        RECT  3.15 0.56 3.31 1.12 ;
        RECT  2.43 0.96 3.31 1.12 ;
        RECT  2.43 0.96 2.71 1.24 ;
        RECT  2.55 0.96 2.71 2.20 ;
        RECT  2.43 1.92 2.71 2.20 ;
        RECT  2.43 2.04 3.31 2.20 ;
        RECT  3.15 2.04 3.31 2.64 ;
        RECT  3.15 2.48 4.35 2.64 ;
        RECT  4.07 2.48 4.35 2.76 ;
        RECT  5.67 0.88 5.95 1.16 ;
        RECT  5.67 0.88 5.83 2.12 ;
        RECT  5.45 1.84 5.83 2.12 ;
        RECT  6.15 1.84 6.43 2.12 ;
        RECT  5.45 1.96 6.43 2.12 ;
        RECT  6.85 0.44 7.13 0.72 ;
        RECT  6.31 0.56 7.13 0.72 ;
        RECT  6.19 0.88 6.47 1.16 ;
        RECT  6.31 0.56 6.47 1.68 ;
        RECT  6.31 1.52 6.75 1.68 ;
        RECT  6.59 1.52 6.75 2.12 ;
        RECT  6.59 1.84 6.95 2.12 ;
        RECT  4.63 0.87 4.91 1.15 ;
        RECT  4.07 0.99 4.91 1.15 ;
        RECT  4.07 0.96 4.35 1.24 ;
        RECT  4.19 0.96 4.35 2.12 ;
        RECT  4.19 1.84 4.47 2.12 ;
        RECT  4.19 1.96 4.77 2.12 ;
        RECT  4.61 1.96 4.77 2.76 ;
        RECT  7.95 2.42 8.23 2.76 ;
        RECT  4.61 2.60 8.23 2.76 ;
        RECT  8.15 0.50 8.43 0.78 ;
        RECT  6.71 0.88 6.99 1.20 ;
        RECT  7.33 0.92 7.61 1.20 ;
        RECT  8.15 0.50 8.31 1.20 ;
        RECT  6.71 1.04 8.31 1.20 ;
        RECT  7.11 1.04 7.27 2.12 ;
        RECT  7.11 1.84 7.47 2.12 ;
        RECT  5.13 0.87 5.43 1.15 ;
        RECT  8.81 0.92 9.09 1.20 ;
        RECT  7.63 1.52 8.97 1.68 ;
        RECT  8.81 0.92 8.97 2.12 ;
        RECT  5.01 1.84 5.29 2.12 ;
        RECT  8.71 1.84 8.99 2.12 ;
        RECT  5.13 0.87 5.29 2.44 ;
        RECT  7.63 1.52 7.79 2.44 ;
        RECT  5.13 2.28 7.79 2.44 ;
        RECT  9.37 0.88 9.65 1.16 ;
        RECT  9.37 1.00 9.91 1.16 ;
        RECT  9.75 1.46 10.75 1.62 ;
        RECT  10.47 1.40 10.75 1.68 ;
        RECT  9.75 1.00 9.91 2.12 ;
        RECT  9.75 1.84 10.03 2.12 ;
        RECT  10.79 0.88 11.07 1.16 ;
        RECT  10.79 1.84 11.07 2.12 ;
        RECT  10.91 0.88 11.07 2.76 ;
        RECT  10.82 2.48 11.10 2.76 ;
        RECT  13.17 0.84 13.45 1.24 ;
        RECT  13.03 1.46 13.33 1.74 ;
        RECT  13.17 0.84 13.33 2.30 ;
        RECT  13.17 1.90 13.45 2.30 ;
    END
END DFFDRHZSP2V1_0

MACRO DFFDRHZSP1V1_0
    CLASS CORE ;
    FOREIGN DFFDRHZSP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.76 2.28 9.14 2.56 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.22 1.40 3.54 1.76 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.20  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.83  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.81 1.19 2.25 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  0.91 0.81 1.19 1.09 ;
        END
    END D
    PIN QZ
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 25.91  LAYER ME1  ;
        ANTENNADIFFAREA 10.52  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.64  LAYER ME1  ;
        ANTENNAMAXAREACAR 40.59  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.73 1.90 13.01 2.18 ;
        RECT  12.73 0.88 13.01 1.16 ;
        RECT  12.73 0.88 12.89 2.18 ;
        RECT  12.46 1.46 12.89 1.74 ;
        END
    END QZ
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 25.91  LAYER ME1  ;
        ANTENNADIFFAREA 10.52  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.64  LAYER ME1  ;
        ANTENNAMAXAREACAR 40.59  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.31 1.90 11.59 2.18 ;
        RECT  11.31 0.88 11.59 1.16 ;
        RECT  11.31 0.88 11.54 2.18 ;
        RECT  11.26 1.46 11.54 1.74 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.10  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.55 1.46 13.95 1.74 ;
        END
    END E
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END SEL
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.87  LAYER ME1  ;
        ANTENNADIFFAREA 0.60  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 12.90  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.06 1.46 2.34 1.74 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.81 2.23 2.25 ;
        RECT  1.95 0.81 2.23 1.09 ;
        END
    END TD
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 14.40 3.48 ;
        RECT  13.79 2.88 14.22 3.48 ;
        RECT  13.73 1.90 14.01 2.18 ;
        RECT  13.79 1.90 13.95 3.48 ;
        RECT  11.83 1.90 12.11 2.18 ;
        RECT  11.89 1.90 12.05 3.48 ;
        RECT  10.27 1.84 10.55 2.12 ;
        RECT  10.33 1.84 10.49 3.48 ;
        RECT  9.43 1.84 9.59 3.48 ;
        RECT  9.23 1.84 9.59 2.12 ;
        RECT  8.39 1.84 8.55 3.48 ;
        RECT  8.19 1.84 8.55 2.12 ;
        RECT  2.71 2.52 2.99 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 14.40 0.28 ;
        RECT  13.78 -0.28 14.22 0.32 ;
        RECT  13.73 0.88 14.01 1.16 ;
        RECT  13.78 -0.28 13.94 1.16 ;
        RECT  11.83 0.88 12.11 1.16 ;
        RECT  11.89 -0.28 12.05 1.16 ;
        RECT  10.27 0.88 10.55 1.16 ;
        RECT  10.33 -0.28 10.49 1.16 ;
        RECT  7.29 -0.28 7.57 0.72 ;
        RECT  2.71 -0.28 2.99 0.68 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  1.55 1.97 1.71 2.57 ;
        RECT  1.55 2.41 2.37 2.57 ;
        RECT  2.09 2.41 2.37 2.69 ;
        RECT  3.47 0.96 3.86 1.24 ;
        RECT  3.70 1.46 4.02 1.74 ;
        RECT  3.70 0.96 3.86 2.20 ;
        RECT  3.47 1.92 3.86 2.20 ;
        RECT  4.07 0.44 4.35 0.72 ;
        RECT  3.15 0.56 4.35 0.72 ;
        RECT  3.15 0.56 3.31 1.12 ;
        RECT  2.43 0.96 3.31 1.12 ;
        RECT  2.43 0.96 2.71 1.24 ;
        RECT  2.55 0.96 2.71 2.20 ;
        RECT  2.43 1.92 2.71 2.20 ;
        RECT  2.43 2.04 3.31 2.20 ;
        RECT  3.15 2.04 3.31 2.64 ;
        RECT  3.15 2.48 4.35 2.64 ;
        RECT  4.07 2.48 4.35 2.76 ;
        RECT  5.67 0.88 5.95 1.16 ;
        RECT  5.67 0.88 5.83 2.12 ;
        RECT  5.45 1.84 5.83 2.12 ;
        RECT  6.15 1.84 6.43 2.12 ;
        RECT  5.45 1.96 6.43 2.12 ;
        RECT  6.85 0.44 7.13 0.72 ;
        RECT  6.31 0.56 7.13 0.72 ;
        RECT  6.19 0.88 6.47 1.16 ;
        RECT  6.31 0.56 6.47 1.68 ;
        RECT  6.31 1.52 6.75 1.68 ;
        RECT  6.59 1.52 6.75 2.12 ;
        RECT  6.59 1.84 6.95 2.12 ;
        RECT  4.63 0.87 4.91 1.15 ;
        RECT  4.07 0.99 4.91 1.15 ;
        RECT  4.07 0.96 4.35 1.24 ;
        RECT  4.19 0.96 4.35 2.12 ;
        RECT  4.19 1.84 4.47 2.12 ;
        RECT  4.19 1.96 4.77 2.12 ;
        RECT  4.61 1.96 4.77 2.76 ;
        RECT  7.95 2.42 8.23 2.76 ;
        RECT  4.61 2.60 8.23 2.76 ;
        RECT  8.15 0.50 8.43 0.78 ;
        RECT  6.71 0.88 6.99 1.20 ;
        RECT  7.33 0.92 7.61 1.20 ;
        RECT  8.15 0.50 8.31 1.20 ;
        RECT  6.71 1.04 8.31 1.20 ;
        RECT  7.11 1.04 7.27 2.12 ;
        RECT  7.11 1.84 7.47 2.12 ;
        RECT  5.13 0.87 5.43 1.15 ;
        RECT  8.81 0.92 9.09 1.20 ;
        RECT  7.63 1.52 8.97 1.68 ;
        RECT  8.81 0.92 8.97 2.12 ;
        RECT  5.01 1.84 5.29 2.12 ;
        RECT  8.71 1.84 8.99 2.12 ;
        RECT  5.13 0.87 5.29 2.44 ;
        RECT  7.63 1.52 7.79 2.44 ;
        RECT  5.13 2.28 7.79 2.44 ;
        RECT  9.37 0.88 9.65 1.16 ;
        RECT  9.37 1.00 9.91 1.16 ;
        RECT  9.75 1.46 10.75 1.62 ;
        RECT  10.47 1.40 10.75 1.68 ;
        RECT  9.75 1.00 9.91 2.12 ;
        RECT  9.75 1.84 10.03 2.12 ;
        RECT  10.79 0.88 11.07 1.16 ;
        RECT  10.79 1.84 11.07 2.12 ;
        RECT  10.91 0.88 11.07 2.76 ;
        RECT  10.82 2.48 11.10 2.76 ;
        RECT  13.21 0.88 13.49 1.16 ;
        RECT  13.07 1.46 13.37 1.74 ;
        RECT  13.21 0.88 13.37 2.18 ;
        RECT  13.21 1.90 13.49 2.18 ;
    END
END DFFDRHZSP1V1_0

MACRO DFFDRHSP8V1_0
    CLASS CORE ;
    FOREIGN DFFDRHSP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.42 2.28 6.80 2.56 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.88 1.40 1.20 1.76 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.40 0.72 1.76 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 30.10  LAYER ME1  ;
        ANTENNADIFFAREA 15.21  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.41  LAYER ME1  ;
        ANTENNAMAXAREACAR 21.33  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.50 1.90 10.78 2.50 ;
        RECT  10.50 0.64 10.78 1.24 ;
        RECT  10.50 0.64 10.66 2.50 ;
        RECT  9.26 1.52 10.66 1.68 ;
        RECT  9.46 1.90 9.74 2.50 ;
        RECT  9.46 0.64 9.74 1.24 ;
        RECT  9.46 0.64 9.62 2.50 ;
        RECT  9.26 1.46 9.62 1.74 ;
        END
    END Q
    PIN QZ
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 30.10  LAYER ME1  ;
        ANTENNADIFFAREA 14.99  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.41  LAYER ME1  ;
        ANTENNAMAXAREACAR 21.33  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.10 1.90 13.38 2.18 ;
        RECT  13.10 0.96 13.38 1.24 ;
        RECT  13.10 0.96 13.26 2.18 ;
        RECT  12.06 1.52 13.26 1.68 ;
        RECT  12.06 0.96 12.34 2.18 ;
        END
    END QZ
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.43  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.44 1.46 14.84 1.74 ;
        END
    END E
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 15.20 0.28 ;
        RECT  14.68 -0.28 15.02 0.32 ;
        RECT  14.62 0.64 14.90 1.24 ;
        RECT  14.68 -0.28 14.84 1.24 ;
        RECT  11.02 0.64 11.30 1.24 ;
        RECT  11.08 -0.28 11.24 1.24 ;
        RECT  9.98 0.64 10.26 1.24 ;
        RECT  10.04 -0.28 10.20 1.24 ;
        RECT  8.94 0.64 9.22 1.24 ;
        RECT  9.00 -0.28 9.16 1.24 ;
        RECT  7.94 0.88 8.22 1.16 ;
        RECT  8.00 -0.28 8.16 1.16 ;
        RECT  4.96 -0.28 5.24 0.72 ;
        RECT  0.38 -0.28 0.66 0.68 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 15.20 3.48 ;
        RECT  14.68 2.88 15.02 3.48 ;
        RECT  14.62 1.90 14.90 2.50 ;
        RECT  14.68 1.90 14.84 3.48 ;
        RECT  11.02 1.90 11.30 2.50 ;
        RECT  11.08 1.90 11.24 3.48 ;
        RECT  9.98 1.90 10.26 2.50 ;
        RECT  10.04 1.90 10.20 3.48 ;
        RECT  8.94 1.90 9.22 2.50 ;
        RECT  9.00 1.90 9.16 3.48 ;
        RECT  7.94 1.84 8.22 2.12 ;
        RECT  8.00 1.84 8.16 3.48 ;
        RECT  7.10 1.84 7.26 3.48 ;
        RECT  6.90 1.84 7.26 2.12 ;
        RECT  6.06 1.84 6.22 3.48 ;
        RECT  5.86 1.84 6.22 2.12 ;
        RECT  0.38 2.48 0.66 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  1.14 0.96 1.52 1.24 ;
        RECT  1.36 1.46 1.64 1.74 ;
        RECT  1.36 0.96 1.52 2.20 ;
        RECT  1.14 1.92 1.52 2.20 ;
        RECT  1.74 0.44 2.02 0.72 ;
        RECT  0.82 0.56 2.02 0.72 ;
        RECT  0.82 0.56 0.98 1.12 ;
        RECT  0.08 0.96 0.98 1.12 ;
        RECT  0.08 0.96 0.38 1.24 ;
        RECT  0.08 0.96 0.24 2.20 ;
        RECT  0.08 1.92 0.38 2.20 ;
        RECT  0.08 2.04 0.98 2.20 ;
        RECT  0.82 2.04 0.98 2.64 ;
        RECT  0.82 2.48 2.02 2.64 ;
        RECT  1.74 2.48 2.02 2.76 ;
        RECT  3.34 0.88 3.62 1.16 ;
        RECT  3.34 0.88 3.50 2.12 ;
        RECT  3.12 1.84 3.50 2.12 ;
        RECT  3.82 1.84 4.10 2.12 ;
        RECT  3.12 1.96 4.10 2.12 ;
        RECT  4.52 0.44 4.80 0.72 ;
        RECT  3.98 0.56 4.80 0.72 ;
        RECT  3.86 0.88 4.14 1.16 ;
        RECT  3.98 0.56 4.14 1.68 ;
        RECT  3.98 1.52 4.42 1.68 ;
        RECT  4.26 1.52 4.42 2.12 ;
        RECT  4.26 1.84 4.62 2.12 ;
        RECT  2.30 0.87 2.58 1.15 ;
        RECT  1.74 0.99 2.58 1.15 ;
        RECT  1.74 0.96 2.02 1.24 ;
        RECT  1.86 0.96 2.02 2.12 ;
        RECT  1.86 1.84 2.14 2.12 ;
        RECT  1.86 1.96 2.44 2.12 ;
        RECT  2.28 1.96 2.44 2.76 ;
        RECT  5.62 2.42 5.90 2.76 ;
        RECT  2.28 2.60 5.90 2.76 ;
        RECT  5.82 0.50 6.10 0.78 ;
        RECT  4.38 0.88 4.66 1.20 ;
        RECT  5.00 0.92 5.28 1.20 ;
        RECT  5.82 0.50 5.98 1.20 ;
        RECT  4.38 1.04 5.98 1.20 ;
        RECT  4.78 1.04 4.94 2.12 ;
        RECT  4.78 1.84 5.14 2.12 ;
        RECT  2.80 0.87 3.10 1.15 ;
        RECT  6.48 0.92 6.76 1.20 ;
        RECT  5.30 1.52 6.64 1.68 ;
        RECT  6.48 0.92 6.64 2.12 ;
        RECT  2.68 1.84 2.96 2.12 ;
        RECT  6.38 1.84 6.66 2.12 ;
        RECT  2.80 0.87 2.96 2.44 ;
        RECT  5.30 1.52 5.46 2.44 ;
        RECT  2.80 2.28 5.46 2.44 ;
        RECT  7.04 0.88 7.32 1.16 ;
        RECT  7.04 1.00 7.58 1.16 ;
        RECT  7.42 1.46 8.42 1.62 ;
        RECT  8.14 1.40 8.42 1.68 ;
        RECT  7.42 1.00 7.58 2.12 ;
        RECT  7.42 1.84 7.70 2.12 ;
        RECT  8.46 0.88 8.74 1.16 ;
        RECT  8.46 1.84 8.74 2.12 ;
        RECT  8.58 0.88 8.74 2.76 ;
        RECT  8.49 2.48 8.77 2.76 ;
        RECT  11.54 1.90 11.82 2.50 ;
        RECT  12.58 1.90 12.86 2.50 ;
        RECT  13.62 1.90 13.90 2.50 ;
        RECT  11.54 2.34 13.90 2.50 ;
        RECT  11.54 0.64 13.90 0.80 ;
        RECT  11.54 0.64 11.82 1.24 ;
        RECT  12.58 0.64 12.86 1.24 ;
        RECT  13.62 0.64 13.90 1.24 ;
        RECT  14.10 0.64 14.38 1.24 ;
        RECT  13.96 1.46 14.26 1.74 ;
        RECT  14.10 0.64 14.26 2.50 ;
        RECT  14.10 1.90 14.38 2.50 ;
    END
END DFFDRHSP8V1_0

MACRO DFFDRHSP4V1_0
    CLASS CORE ;
    FOREIGN DFFDRHSP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 13.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.26  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.36 1.46 12.76 1.74 ;
        END
    END E
    PIN QZ
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 25.44  LAYER ME1  ;
        ANTENNADIFFAREA 12.29  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.98  LAYER ME1  ;
        ANTENNAMAXAREACAR 25.98  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.02 1.90 11.30 2.18 ;
        RECT  11.02 0.96 11.30 1.24 ;
        RECT  11.02 0.96 11.18 2.18 ;
        RECT  10.86 1.46 11.18 1.74 ;
        END
    END QZ
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 25.74  LAYER ME1  ;
        ANTENNADIFFAREA 12.27  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.98  LAYER ME1  ;
        ANTENNAMAXAREACAR 26.29  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.46 1.90 9.74 2.50 ;
        RECT  9.46 0.64 9.74 1.24 ;
        RECT  9.46 0.64 9.62 2.50 ;
        RECT  9.26 1.46 9.62 1.74 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.40 0.72 1.76 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.88 1.40 1.20 1.76 ;
        END
    END CK
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.42 2.28 6.80 2.56 ;
        END
    END RB
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 13.20 0.28 ;
        RECT  12.60 -0.28 13.02 0.32 ;
        RECT  12.54 0.74 12.82 1.24 ;
        RECT  12.60 -0.28 12.76 1.24 ;
        RECT  9.98 0.64 10.26 1.24 ;
        RECT  10.04 -0.28 10.20 1.24 ;
        RECT  8.94 0.64 9.22 1.24 ;
        RECT  9.00 -0.28 9.16 1.24 ;
        RECT  7.94 0.88 8.22 1.16 ;
        RECT  8.00 -0.28 8.16 1.16 ;
        RECT  4.96 -0.28 5.24 0.72 ;
        RECT  0.38 -0.28 0.66 0.68 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 13.20 3.48 ;
        RECT  12.60 2.88 13.02 3.48 ;
        RECT  12.54 1.90 12.82 2.40 ;
        RECT  12.60 1.90 12.76 3.48 ;
        RECT  9.98 1.90 10.26 2.50 ;
        RECT  10.04 1.90 10.20 3.48 ;
        RECT  8.94 1.90 9.22 2.50 ;
        RECT  9.00 1.90 9.16 3.48 ;
        RECT  7.94 1.84 8.22 2.12 ;
        RECT  8.00 1.84 8.16 3.48 ;
        RECT  7.10 1.84 7.26 3.48 ;
        RECT  6.90 1.84 7.26 2.12 ;
        RECT  6.06 1.84 6.22 3.48 ;
        RECT  5.86 1.84 6.22 2.12 ;
        RECT  0.38 2.48 0.66 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  1.14 0.96 1.52 1.24 ;
        RECT  1.36 1.46 1.64 1.74 ;
        RECT  1.36 0.96 1.52 2.20 ;
        RECT  1.14 1.92 1.52 2.20 ;
        RECT  1.74 0.44 2.02 0.72 ;
        RECT  0.82 0.56 2.02 0.72 ;
        RECT  0.82 0.56 0.98 1.12 ;
        RECT  0.08 0.96 0.98 1.12 ;
        RECT  0.08 0.96 0.38 1.24 ;
        RECT  0.08 0.96 0.24 2.20 ;
        RECT  0.08 1.92 0.38 2.20 ;
        RECT  0.08 2.04 0.98 2.20 ;
        RECT  0.82 2.04 0.98 2.64 ;
        RECT  0.82 2.48 2.02 2.64 ;
        RECT  1.74 2.48 2.02 2.76 ;
        RECT  3.34 0.88 3.62 1.16 ;
        RECT  3.34 0.88 3.50 2.12 ;
        RECT  3.12 1.84 3.50 2.12 ;
        RECT  3.82 1.84 4.10 2.12 ;
        RECT  3.12 1.96 4.10 2.12 ;
        RECT  4.52 0.44 4.80 0.72 ;
        RECT  3.98 0.56 4.80 0.72 ;
        RECT  3.86 0.88 4.14 1.16 ;
        RECT  3.98 0.56 4.14 1.68 ;
        RECT  3.98 1.52 4.42 1.68 ;
        RECT  4.26 1.52 4.42 2.12 ;
        RECT  4.26 1.84 4.62 2.12 ;
        RECT  2.30 0.87 2.58 1.15 ;
        RECT  1.74 0.99 2.58 1.15 ;
        RECT  1.74 0.96 2.02 1.24 ;
        RECT  1.86 0.96 2.02 2.12 ;
        RECT  1.86 1.84 2.14 2.12 ;
        RECT  1.86 1.96 2.44 2.12 ;
        RECT  2.28 1.96 2.44 2.76 ;
        RECT  5.62 2.42 5.90 2.76 ;
        RECT  2.28 2.60 5.90 2.76 ;
        RECT  5.82 0.50 6.10 0.78 ;
        RECT  4.38 0.88 4.66 1.20 ;
        RECT  5.00 0.92 5.28 1.20 ;
        RECT  5.82 0.50 5.98 1.20 ;
        RECT  4.38 1.04 5.98 1.20 ;
        RECT  4.78 1.04 4.94 2.12 ;
        RECT  4.78 1.84 5.14 2.12 ;
        RECT  2.80 0.87 3.10 1.15 ;
        RECT  6.48 0.92 6.76 1.20 ;
        RECT  5.30 1.52 6.64 1.68 ;
        RECT  6.48 0.92 6.64 2.12 ;
        RECT  2.68 1.84 2.96 2.12 ;
        RECT  6.38 1.84 6.66 2.12 ;
        RECT  2.80 0.87 2.96 2.44 ;
        RECT  5.30 1.52 5.46 2.44 ;
        RECT  2.80 2.28 5.46 2.44 ;
        RECT  7.04 0.88 7.32 1.16 ;
        RECT  7.04 1.00 7.58 1.16 ;
        RECT  7.42 1.46 8.42 1.62 ;
        RECT  8.14 1.40 8.42 1.68 ;
        RECT  7.42 1.00 7.58 2.12 ;
        RECT  7.42 1.84 7.70 2.12 ;
        RECT  8.46 0.88 8.74 1.16 ;
        RECT  8.46 1.84 8.74 2.12 ;
        RECT  8.58 0.88 8.74 2.76 ;
        RECT  8.49 2.48 8.77 2.76 ;
        RECT  10.50 1.90 10.78 2.50 ;
        RECT  11.54 1.90 11.82 2.50 ;
        RECT  10.50 2.34 11.82 2.50 ;
        RECT  10.50 0.64 11.82 0.80 ;
        RECT  10.50 0.64 10.78 1.24 ;
        RECT  11.54 0.64 11.82 1.24 ;
        RECT  12.02 0.74 12.30 1.24 ;
        RECT  11.88 1.46 12.18 1.74 ;
        RECT  12.02 0.74 12.18 2.40 ;
        RECT  12.02 1.90 12.30 2.40 ;
    END
END DFFDRHSP4V1_0

MACRO DFFDRHSP2V1_0
    CLASS CORE ;
    FOREIGN DFFDRHSP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.42 2.28 6.80 2.56 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.88 1.40 1.20 1.76 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.40 0.72 1.76 ;
        END
    END D
    PIN QZ
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 23.19  LAYER ME1  ;
        ANTENNADIFFAREA 10.39  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.76  LAYER ME1  ;
        ANTENNAMAXAREACAR 30.39  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.36 1.90 10.64 2.50 ;
        RECT  10.36 0.64 10.64 1.24 ;
        RECT  10.36 0.64 10.52 2.50 ;
        RECT  10.06 1.46 10.52 1.74 ;
        END
    END QZ
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 23.19  LAYER ME1  ;
        ANTENNADIFFAREA 10.39  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.76  LAYER ME1  ;
        ANTENNAMAXAREACAR 30.39  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.06 1.46 9.54 1.74 ;
        RECT  8.94 1.90 9.22 2.50 ;
        RECT  9.06 0.64 9.22 2.50 ;
        RECT  8.94 0.64 9.22 1.24 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.17  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.16 1.46 11.56 1.74 ;
        END
    END E
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 12.00 3.48 ;
        RECT  11.42 2.88 11.82 3.48 ;
        RECT  11.36 1.90 11.64 2.30 ;
        RECT  11.42 1.90 11.58 3.48 ;
        RECT  9.46 1.90 9.74 2.50 ;
        RECT  9.52 1.90 9.68 3.48 ;
        RECT  7.94 1.84 8.22 2.12 ;
        RECT  8.00 1.84 8.16 3.48 ;
        RECT  7.10 1.84 7.26 3.48 ;
        RECT  6.90 1.84 7.26 2.12 ;
        RECT  6.06 1.84 6.22 3.48 ;
        RECT  5.86 1.84 6.22 2.12 ;
        RECT  0.38 2.48 0.66 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 12.00 0.28 ;
        RECT  11.42 -0.28 11.82 0.32 ;
        RECT  11.36 0.84 11.64 1.24 ;
        RECT  11.42 -0.28 11.58 1.24 ;
        RECT  9.46 0.64 9.74 1.24 ;
        RECT  9.52 -0.28 9.68 1.24 ;
        RECT  7.94 0.88 8.22 1.16 ;
        RECT  8.00 -0.28 8.16 1.16 ;
        RECT  4.96 -0.28 5.24 0.72 ;
        RECT  0.38 -0.28 0.66 0.68 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  1.14 0.96 1.52 1.24 ;
        RECT  1.36 1.46 1.64 1.74 ;
        RECT  1.36 0.96 1.52 2.20 ;
        RECT  1.14 1.92 1.52 2.20 ;
        RECT  1.74 0.44 2.02 0.72 ;
        RECT  0.82 0.56 2.02 0.72 ;
        RECT  0.82 0.56 0.98 1.12 ;
        RECT  0.08 0.96 0.98 1.12 ;
        RECT  0.08 0.96 0.38 1.24 ;
        RECT  0.08 0.96 0.24 2.20 ;
        RECT  0.08 1.92 0.38 2.20 ;
        RECT  0.08 2.04 0.98 2.20 ;
        RECT  0.82 2.04 0.98 2.64 ;
        RECT  0.82 2.48 2.02 2.64 ;
        RECT  1.74 2.48 2.02 2.76 ;
        RECT  3.34 0.88 3.62 1.16 ;
        RECT  3.34 0.88 3.50 2.12 ;
        RECT  3.12 1.84 3.50 2.12 ;
        RECT  3.82 1.84 4.10 2.12 ;
        RECT  3.12 1.96 4.10 2.12 ;
        RECT  4.52 0.44 4.80 0.72 ;
        RECT  3.98 0.56 4.80 0.72 ;
        RECT  3.86 0.88 4.14 1.16 ;
        RECT  3.98 0.56 4.14 1.68 ;
        RECT  3.98 1.52 4.42 1.68 ;
        RECT  4.26 1.52 4.42 2.12 ;
        RECT  4.26 1.84 4.62 2.12 ;
        RECT  2.30 0.87 2.58 1.15 ;
        RECT  1.74 0.99 2.58 1.15 ;
        RECT  1.74 0.96 2.02 1.24 ;
        RECT  1.86 0.96 2.02 2.12 ;
        RECT  1.86 1.84 2.14 2.12 ;
        RECT  1.86 1.96 2.44 2.12 ;
        RECT  2.28 1.96 2.44 2.76 ;
        RECT  5.62 2.42 5.90 2.76 ;
        RECT  2.28 2.60 5.90 2.76 ;
        RECT  5.82 0.50 6.10 0.78 ;
        RECT  4.38 0.88 4.66 1.20 ;
        RECT  5.00 0.92 5.28 1.20 ;
        RECT  5.82 0.50 5.98 1.20 ;
        RECT  4.38 1.04 5.98 1.20 ;
        RECT  4.78 1.04 4.94 2.12 ;
        RECT  4.78 1.84 5.14 2.12 ;
        RECT  2.80 0.87 3.10 1.15 ;
        RECT  6.48 0.92 6.76 1.20 ;
        RECT  5.30 1.52 6.64 1.68 ;
        RECT  6.48 0.92 6.64 2.12 ;
        RECT  2.68 1.84 2.96 2.12 ;
        RECT  6.38 1.84 6.66 2.12 ;
        RECT  2.80 0.87 2.96 2.44 ;
        RECT  5.30 1.52 5.46 2.44 ;
        RECT  2.80 2.28 5.46 2.44 ;
        RECT  7.04 0.88 7.32 1.16 ;
        RECT  7.04 1.00 7.58 1.16 ;
        RECT  7.42 1.46 8.42 1.62 ;
        RECT  8.14 1.40 8.42 1.68 ;
        RECT  7.42 1.00 7.58 2.12 ;
        RECT  7.42 1.84 7.70 2.12 ;
        RECT  8.46 0.88 8.74 1.16 ;
        RECT  8.46 1.84 8.74 2.12 ;
        RECT  8.58 0.88 8.74 2.76 ;
        RECT  8.49 2.48 8.77 2.76 ;
        RECT  10.84 0.84 11.12 1.24 ;
        RECT  10.70 1.46 11.00 1.74 ;
        RECT  10.84 0.84 11.00 2.30 ;
        RECT  10.84 1.90 11.12 2.30 ;
    END
END DFFDRHSP2V1_0

MACRO DFFDRHSP1V1_0
    CLASS CORE ;
    FOREIGN DFFDRHSP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 22.67  LAYER ME1  ;
        ANTENNADIFFAREA 9.37  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER ME1  ;
        ANTENNAMAXAREACAR 39.69  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.10 1.46 9.54 1.74 ;
        RECT  8.98 1.90 9.26 2.18 ;
        RECT  9.10 0.88 9.26 2.18 ;
        RECT  8.98 0.88 9.26 1.16 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.10  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.22 1.46 11.62 1.74 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.40 0.72 1.76 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.88 1.40 1.20 1.76 ;
        END
    END CK
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.42 2.28 6.80 2.56 ;
        END
    END RB
    PIN QZ
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 22.67  LAYER ME1  ;
        ANTENNADIFFAREA 9.37  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER ME1  ;
        ANTENNAMAXAREACAR 39.69  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.40 1.90 10.68 2.18 ;
        RECT  10.40 0.88 10.68 1.16 ;
        RECT  10.40 0.88 10.56 2.18 ;
        RECT  10.06 1.46 10.56 1.74 ;
        END
    END QZ
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 12.00 0.28 ;
        RECT  11.45 -0.28 11.82 0.32 ;
        RECT  11.40 0.88 11.68 1.16 ;
        RECT  11.45 -0.28 11.61 1.16 ;
        RECT  9.50 0.88 9.78 1.16 ;
        RECT  9.56 -0.28 9.72 1.16 ;
        RECT  7.94 0.88 8.22 1.16 ;
        RECT  8.00 -0.28 8.16 1.16 ;
        RECT  4.96 -0.28 5.24 0.72 ;
        RECT  0.38 -0.28 0.66 0.68 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 12.00 3.48 ;
        RECT  11.46 2.88 11.82 3.48 ;
        RECT  11.40 1.90 11.68 2.18 ;
        RECT  11.46 1.90 11.62 3.48 ;
        RECT  9.50 1.90 9.78 2.18 ;
        RECT  9.56 1.90 9.72 3.48 ;
        RECT  7.94 1.84 8.22 2.12 ;
        RECT  8.00 1.84 8.16 3.48 ;
        RECT  7.10 1.84 7.26 3.48 ;
        RECT  6.90 1.84 7.26 2.12 ;
        RECT  6.06 1.84 6.22 3.48 ;
        RECT  5.86 1.84 6.22 2.12 ;
        RECT  0.38 2.48 0.66 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  1.14 0.96 1.52 1.24 ;
        RECT  1.36 1.46 1.64 1.74 ;
        RECT  1.36 0.96 1.52 2.20 ;
        RECT  1.14 1.92 1.52 2.20 ;
        RECT  1.74 0.44 2.02 0.72 ;
        RECT  0.82 0.56 2.02 0.72 ;
        RECT  0.82 0.56 0.98 1.12 ;
        RECT  0.08 0.96 0.98 1.12 ;
        RECT  0.08 0.96 0.38 1.24 ;
        RECT  0.08 0.96 0.24 2.20 ;
        RECT  0.08 1.92 0.38 2.20 ;
        RECT  0.08 2.04 0.98 2.20 ;
        RECT  0.82 2.04 0.98 2.64 ;
        RECT  0.82 2.48 2.02 2.64 ;
        RECT  1.74 2.48 2.02 2.76 ;
        RECT  3.34 0.88 3.62 1.16 ;
        RECT  3.34 0.88 3.50 2.12 ;
        RECT  3.12 1.84 3.50 2.12 ;
        RECT  3.82 1.84 4.10 2.12 ;
        RECT  3.12 1.96 4.10 2.12 ;
        RECT  4.52 0.44 4.80 0.72 ;
        RECT  3.98 0.56 4.80 0.72 ;
        RECT  3.86 0.88 4.14 1.16 ;
        RECT  3.98 0.56 4.14 1.68 ;
        RECT  3.98 1.52 4.42 1.68 ;
        RECT  4.26 1.52 4.42 2.12 ;
        RECT  4.26 1.84 4.62 2.12 ;
        RECT  2.30 0.87 2.58 1.15 ;
        RECT  1.74 0.99 2.58 1.15 ;
        RECT  1.74 0.96 2.02 1.24 ;
        RECT  1.86 0.96 2.02 2.12 ;
        RECT  1.86 1.84 2.14 2.12 ;
        RECT  1.86 1.96 2.44 2.12 ;
        RECT  2.28 1.96 2.44 2.76 ;
        RECT  5.62 2.42 5.90 2.76 ;
        RECT  2.28 2.60 5.90 2.76 ;
        RECT  5.82 0.50 6.10 0.78 ;
        RECT  4.38 0.88 4.66 1.20 ;
        RECT  5.00 0.92 5.28 1.20 ;
        RECT  5.82 0.50 5.98 1.20 ;
        RECT  4.38 1.04 5.98 1.20 ;
        RECT  4.78 1.04 4.94 2.12 ;
        RECT  4.78 1.84 5.14 2.12 ;
        RECT  2.80 0.87 3.10 1.15 ;
        RECT  6.48 0.92 6.76 1.20 ;
        RECT  5.30 1.52 6.64 1.68 ;
        RECT  6.48 0.92 6.64 2.12 ;
        RECT  2.68 1.84 2.96 2.12 ;
        RECT  6.38 1.84 6.66 2.12 ;
        RECT  2.80 0.87 2.96 2.44 ;
        RECT  5.30 1.52 5.46 2.44 ;
        RECT  2.80 2.28 5.46 2.44 ;
        RECT  7.04 0.88 7.32 1.16 ;
        RECT  7.04 1.00 7.58 1.16 ;
        RECT  7.42 1.46 8.42 1.62 ;
        RECT  8.14 1.40 8.42 1.68 ;
        RECT  7.42 1.00 7.58 2.12 ;
        RECT  7.42 1.84 7.70 2.12 ;
        RECT  8.46 0.88 8.74 1.16 ;
        RECT  8.46 1.84 8.74 2.12 ;
        RECT  8.58 0.88 8.74 2.76 ;
        RECT  8.49 2.48 8.77 2.76 ;
        RECT  10.88 0.88 11.16 1.16 ;
        RECT  10.74 1.46 11.04 1.74 ;
        RECT  10.88 0.88 11.04 2.18 ;
        RECT  10.88 1.90 11.16 2.18 ;
    END
END DFFDRHSP1V1_0

MACRO DFFDRBZSP8V1_0
    CLASS CORE ;
    FOREIGN DFFDRBZSP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 27.30  LAYER ME1  ;
        ANTENNADIFFAREA 13.99  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.62  LAYER ME1  ;
        ANTENNAMAXAREACAR 16.83  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.78 1.90 14.06 2.18 ;
        RECT  13.78 0.96 14.06 1.24 ;
        RECT  13.78 0.96 13.94 2.18 ;
        RECT  12.86 1.52 13.94 1.68 ;
        RECT  12.86 1.46 13.14 1.74 ;
        RECT  12.74 1.90 13.02 2.18 ;
        RECT  12.86 0.96 13.02 2.18 ;
        RECT  12.74 0.96 13.02 1.24 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 27.30  LAYER ME1  ;
        ANTENNADIFFAREA 13.99  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.62  LAYER ME1  ;
        ANTENNAMAXAREACAR 16.83  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.70 1.90 11.98 2.18 ;
        RECT  11.70 0.96 11.98 1.24 ;
        RECT  11.70 0.96 11.86 2.18 ;
        RECT  10.78 1.52 11.86 1.68 ;
        RECT  10.78 1.46 11.14 1.74 ;
        RECT  10.66 1.90 10.94 2.18 ;
        RECT  10.78 0.96 10.94 2.18 ;
        RECT  10.66 0.96 10.94 1.24 ;
        END
    END QB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.02 1.25 4.30 1.70 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END D
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.42 1.62 1.78 ;
        END
    END SEL
    PIN TD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.62 1.86 3.94 2.14 ;
        RECT  3.62 1.42 3.78 2.14 ;
        RECT  3.42 1.42 3.78 1.70 ;
        END
    END TD
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.36 1.14 1.78 ;
        END
    END RB
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 14.80 0.28 ;
        RECT  14.34 -0.28 14.62 0.32 ;
        RECT  14.30 0.64 14.58 0.92 ;
        RECT  14.36 -0.28 14.52 0.92 ;
        RECT  13.26 0.64 13.54 0.92 ;
        RECT  13.32 -0.28 13.48 0.92 ;
        RECT  12.22 0.64 12.50 0.92 ;
        RECT  12.28 -0.28 12.44 0.92 ;
        RECT  11.18 0.64 11.46 0.92 ;
        RECT  11.24 -0.28 11.40 0.92 ;
        RECT  10.14 0.64 10.42 0.92 ;
        RECT  10.20 -0.28 10.36 0.92 ;
        RECT  9.14 0.96 9.42 1.24 ;
        RECT  9.24 -0.28 9.40 1.24 ;
        RECT  6.40 0.72 6.68 1.00 ;
        RECT  6.46 -0.28 6.62 1.00 ;
        RECT  3.70 0.68 3.98 0.96 ;
        RECT  3.76 -0.28 3.92 0.96 ;
        RECT  1.14 0.70 1.42 0.98 ;
        RECT  1.20 -0.28 1.36 0.98 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 14.80 3.48 ;
        RECT  14.34 2.88 14.62 3.48 ;
        RECT  14.30 2.22 14.58 2.50 ;
        RECT  14.36 2.22 14.52 3.48 ;
        RECT  13.26 2.22 13.54 2.50 ;
        RECT  13.32 2.22 13.48 3.48 ;
        RECT  12.22 2.22 12.50 2.50 ;
        RECT  12.28 2.22 12.44 3.48 ;
        RECT  11.18 2.22 11.46 2.50 ;
        RECT  11.24 2.22 11.40 3.48 ;
        RECT  10.14 1.90 10.42 2.18 ;
        RECT  10.20 1.90 10.36 3.48 ;
        RECT  9.14 2.62 9.42 3.48 ;
        RECT  6.58 1.92 6.86 2.20 ;
        RECT  6.64 1.92 6.80 3.48 ;
        RECT  3.70 2.62 3.98 3.48 ;
        RECT  0.92 2.62 1.20 3.48 ;
        RECT  0.10 1.94 0.38 2.22 ;
        RECT  0.16 1.94 0.32 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  1.66 0.70 1.94 0.98 ;
        RECT  1.78 1.20 2.10 1.48 ;
        RECT  1.78 0.70 1.94 2.22 ;
        RECT  1.66 1.94 1.94 2.22 ;
        RECT  0.10 0.70 0.38 0.98 ;
        RECT  2.14 0.68 2.42 0.96 ;
        RECT  0.10 0.82 0.70 0.98 ;
        RECT  0.54 0.82 0.70 2.22 ;
        RECT  0.54 1.94 0.90 2.22 ;
        RECT  2.26 0.68 2.42 2.14 ;
        RECT  0.54 2.06 1.50 2.22 ;
        RECT  1.34 2.06 1.50 2.54 ;
        RECT  2.14 1.86 2.30 2.54 ;
        RECT  1.34 2.38 2.30 2.54 ;
        RECT  3.10 0.68 3.46 0.96 ;
        RECT  3.10 0.68 3.26 2.14 ;
        RECT  3.10 1.86 3.46 2.14 ;
        RECT  4.22 0.68 4.62 0.96 ;
        RECT  4.46 1.16 4.82 1.44 ;
        RECT  4.46 0.68 4.62 2.14 ;
        RECT  4.22 1.86 4.62 2.14 ;
        RECT  2.66 0.68 2.94 0.96 ;
        RECT  4.78 0.72 5.14 1.00 ;
        RECT  2.72 0.68 2.88 2.14 ;
        RECT  2.66 1.86 2.94 2.14 ;
        RECT  4.98 0.72 5.14 2.20 ;
        RECT  4.78 1.92 5.14 2.20 ;
        RECT  2.78 1.86 2.94 2.46 ;
        RECT  4.78 1.92 4.94 2.46 ;
        RECT  2.78 2.30 4.94 2.46 ;
        RECT  5.86 0.72 6.16 1.00 ;
        RECT  5.86 0.72 6.02 2.20 ;
        RECT  5.82 1.92 6.10 2.20 ;
        RECT  5.30 0.72 5.58 1.00 ;
        RECT  6.66 1.48 6.94 1.76 ;
        RECT  6.26 1.60 6.94 1.76 ;
        RECT  5.36 0.72 5.52 2.20 ;
        RECT  5.30 1.92 5.58 2.20 ;
        RECT  5.42 1.92 5.58 2.52 ;
        RECT  6.26 1.60 6.42 2.52 ;
        RECT  5.42 2.36 6.42 2.52 ;
        RECT  6.92 0.72 7.26 1.00 ;
        RECT  6.18 1.16 7.26 1.32 ;
        RECT  6.18 1.16 6.46 1.44 ;
        RECT  7.10 0.72 7.26 2.20 ;
        RECT  7.10 1.92 7.38 2.20 ;
        RECT  7.60 0.44 9.08 0.60 ;
        RECT  8.80 0.44 9.08 0.80 ;
        RECT  7.48 0.76 7.76 1.04 ;
        RECT  7.60 0.44 7.76 2.20 ;
        RECT  7.60 1.92 7.90 2.20 ;
        RECT  8.62 0.96 8.90 1.24 ;
        RECT  8.62 1.46 9.56 1.62 ;
        RECT  9.28 1.40 9.56 1.68 ;
        RECT  8.62 0.96 8.78 2.12 ;
        RECT  8.62 1.84 8.90 2.12 ;
        RECT  8.00 0.76 8.30 1.04 ;
        RECT  9.66 0.96 9.94 1.24 ;
        RECT  9.66 1.84 9.94 2.12 ;
        RECT  8.14 0.76 8.30 2.20 ;
        RECT  8.26 1.92 8.42 2.44 ;
        RECT  9.75 0.96 9.91 2.70 ;
        RECT  8.26 2.28 9.91 2.44 ;
        RECT  9.75 2.42 10.04 2.70 ;
    END
END DFFDRBZSP8V1_0

MACRO DFFDRBZSP4V1_0
    CLASS CORE ;
    FOREIGN DFFDRBZSP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.36 1.14 1.78 ;
        END
    END RB
    PIN TD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.62 1.86 3.94 2.14 ;
        RECT  3.62 1.42 3.78 2.14 ;
        RECT  3.42 1.42 3.78 1.70 ;
        END
    END TD
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.42 1.62 1.78 ;
        END
    END SEL
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.02 1.25 4.30 1.70 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 23.82  LAYER ME1  ;
        ANTENNADIFFAREA 11.22  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.05  LAYER ME1  ;
        ANTENNAMAXAREACAR 22.76  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.78 1.46 11.14 1.74 ;
        RECT  10.66 1.90 10.94 2.18 ;
        RECT  10.78 0.96 10.94 2.18 ;
        RECT  10.66 0.96 10.94 1.24 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 23.82  LAYER ME1  ;
        ANTENNADIFFAREA 11.22  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.05  LAYER ME1  ;
        ANTENNAMAXAREACAR 22.76  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.70 1.90 11.98 2.18 ;
        RECT  11.70 0.96 11.98 1.24 ;
        RECT  11.70 0.96 11.94 2.18 ;
        RECT  11.66 1.46 11.94 1.74 ;
        END
    END Q
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 12.80 0.28 ;
        RECT  12.28 -0.28 12.62 0.32 ;
        RECT  12.22 0.64 12.50 0.92 ;
        RECT  12.28 -0.28 12.44 0.92 ;
        RECT  11.18 0.64 11.46 0.92 ;
        RECT  11.24 -0.28 11.40 0.92 ;
        RECT  10.14 0.64 10.42 0.92 ;
        RECT  10.20 -0.28 10.36 0.92 ;
        RECT  9.14 0.96 9.42 1.24 ;
        RECT  9.24 -0.28 9.40 1.24 ;
        RECT  6.40 0.72 6.68 1.00 ;
        RECT  6.46 -0.28 6.62 1.00 ;
        RECT  3.70 0.68 3.98 0.96 ;
        RECT  3.76 -0.28 3.92 0.96 ;
        RECT  1.14 0.70 1.42 0.98 ;
        RECT  1.20 -0.28 1.36 0.98 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 12.80 3.48 ;
        RECT  12.28 2.88 12.62 3.48 ;
        RECT  12.22 2.22 12.50 2.50 ;
        RECT  12.28 2.22 12.44 3.48 ;
        RECT  11.18 2.22 11.46 2.50 ;
        RECT  11.24 2.22 11.40 3.48 ;
        RECT  10.14 1.90 10.42 2.18 ;
        RECT  10.20 1.90 10.36 3.48 ;
        RECT  9.14 2.62 9.42 3.48 ;
        RECT  6.58 1.92 6.86 2.20 ;
        RECT  6.64 1.92 6.80 3.48 ;
        RECT  3.70 2.62 3.98 3.48 ;
        RECT  0.92 2.62 1.20 3.48 ;
        RECT  0.10 1.94 0.38 2.22 ;
        RECT  0.16 1.94 0.32 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  1.66 0.70 1.94 0.98 ;
        RECT  1.78 1.20 2.10 1.48 ;
        RECT  1.78 0.70 1.94 2.22 ;
        RECT  1.66 1.94 1.94 2.22 ;
        RECT  0.10 0.70 0.38 0.98 ;
        RECT  2.14 0.68 2.42 0.96 ;
        RECT  0.10 0.82 0.70 0.98 ;
        RECT  0.54 0.82 0.70 2.22 ;
        RECT  0.54 1.94 0.90 2.22 ;
        RECT  2.26 0.68 2.42 2.14 ;
        RECT  0.54 2.06 1.50 2.22 ;
        RECT  1.34 2.06 1.50 2.54 ;
        RECT  2.14 1.86 2.30 2.54 ;
        RECT  1.34 2.38 2.30 2.54 ;
        RECT  3.10 0.68 3.46 0.96 ;
        RECT  3.10 0.68 3.26 2.14 ;
        RECT  3.10 1.86 3.46 2.14 ;
        RECT  4.22 0.68 4.62 0.96 ;
        RECT  4.46 1.16 4.82 1.44 ;
        RECT  4.46 0.68 4.62 2.14 ;
        RECT  4.22 1.86 4.62 2.14 ;
        RECT  2.66 0.68 2.94 0.96 ;
        RECT  4.78 0.72 5.14 1.00 ;
        RECT  2.72 0.68 2.88 2.14 ;
        RECT  2.66 1.86 2.94 2.14 ;
        RECT  4.98 0.72 5.14 2.20 ;
        RECT  4.78 1.92 5.14 2.20 ;
        RECT  2.78 1.86 2.94 2.46 ;
        RECT  4.78 1.92 4.94 2.46 ;
        RECT  2.78 2.30 4.94 2.46 ;
        RECT  5.86 0.72 6.16 1.00 ;
        RECT  5.86 0.72 6.02 2.20 ;
        RECT  5.82 1.92 6.10 2.20 ;
        RECT  5.30 0.72 5.58 1.00 ;
        RECT  6.66 1.48 6.94 1.76 ;
        RECT  6.26 1.60 6.94 1.76 ;
        RECT  5.36 0.72 5.52 2.20 ;
        RECT  5.30 1.92 5.58 2.20 ;
        RECT  5.42 1.92 5.58 2.52 ;
        RECT  6.26 1.60 6.42 2.52 ;
        RECT  5.42 2.36 6.42 2.52 ;
        RECT  6.92 0.72 7.26 1.00 ;
        RECT  6.18 1.16 7.26 1.32 ;
        RECT  6.18 1.16 6.46 1.44 ;
        RECT  7.10 0.72 7.26 2.20 ;
        RECT  7.10 1.92 7.38 2.20 ;
        RECT  7.60 0.44 9.08 0.60 ;
        RECT  8.80 0.44 9.08 0.80 ;
        RECT  7.48 0.76 7.76 1.04 ;
        RECT  7.60 0.44 7.76 2.20 ;
        RECT  7.60 1.92 7.90 2.20 ;
        RECT  8.62 0.96 8.90 1.24 ;
        RECT  8.62 1.46 9.56 1.62 ;
        RECT  9.28 1.40 9.56 1.68 ;
        RECT  8.62 0.96 8.78 2.12 ;
        RECT  8.62 1.84 8.90 2.12 ;
        RECT  8.00 0.76 8.30 1.04 ;
        RECT  9.66 0.96 9.94 1.24 ;
        RECT  9.66 1.84 9.94 2.12 ;
        RECT  8.14 0.76 8.30 2.20 ;
        RECT  8.26 1.92 8.42 2.44 ;
        RECT  9.75 0.96 9.91 2.70 ;
        RECT  8.26 2.28 9.91 2.44 ;
        RECT  9.75 2.42 10.04 2.70 ;
    END
END DFFDRBZSP4V1_0

MACRO DFFDRBZSP2V1_0
    CLASS CORE ;
    FOREIGN DFFDRBZSP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 21.58  LAYER ME1  ;
        ANTENNADIFFAREA 9.85  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.76  LAYER ME1  ;
        ANTENNAMAXAREACAR 28.45  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.26 1.46 11.52 1.74 ;
        RECT  11.18 1.90 11.46 2.18 ;
        RECT  11.26 0.96 11.46 2.18 ;
        RECT  11.18 0.96 11.46 1.24 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 21.88  LAYER ME1  ;
        ANTENNADIFFAREA 9.85  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.76  LAYER ME1  ;
        ANTENNAMAXAREACAR 28.85  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.26 1.46 10.74 1.74 ;
        RECT  10.14 1.90 10.42 2.18 ;
        RECT  10.26 0.96 10.42 2.18 ;
        RECT  10.14 0.96 10.42 1.24 ;
        END
    END QB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.02 1.25 4.30 1.70 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END D
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.42 1.62 1.78 ;
        END
    END SEL
    PIN TD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.62 1.86 3.94 2.14 ;
        RECT  3.62 1.42 3.78 2.14 ;
        RECT  3.42 1.42 3.78 1.70 ;
        END
    END TD
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.36 1.14 1.78 ;
        END
    END RB
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 11.60 3.48 ;
        RECT  11.14 2.88 11.42 3.48 ;
        RECT  10.66 2.22 10.94 2.50 ;
        RECT  10.72 2.22 10.88 3.48 ;
        RECT  9.14 2.62 9.42 3.48 ;
        RECT  6.58 1.92 6.86 2.20 ;
        RECT  6.64 1.92 6.80 3.48 ;
        RECT  3.70 2.62 3.98 3.48 ;
        RECT  0.92 2.62 1.20 3.48 ;
        RECT  0.10 1.94 0.38 2.22 ;
        RECT  0.16 1.94 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 11.60 0.28 ;
        RECT  11.14 -0.28 11.42 0.32 ;
        RECT  10.66 0.64 10.94 0.92 ;
        RECT  10.72 -0.28 10.88 0.92 ;
        RECT  9.14 0.96 9.42 1.24 ;
        RECT  9.24 -0.28 9.40 1.24 ;
        RECT  6.40 0.72 6.68 1.00 ;
        RECT  6.46 -0.28 6.62 1.00 ;
        RECT  3.70 0.68 3.98 0.96 ;
        RECT  3.76 -0.28 3.92 0.96 ;
        RECT  1.14 0.70 1.42 0.98 ;
        RECT  1.20 -0.28 1.36 0.98 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  1.66 0.70 1.94 0.98 ;
        RECT  1.78 1.20 2.10 1.48 ;
        RECT  1.78 0.70 1.94 2.22 ;
        RECT  1.66 1.94 1.94 2.22 ;
        RECT  0.10 0.70 0.38 0.98 ;
        RECT  2.14 0.68 2.42 0.96 ;
        RECT  0.10 0.82 0.70 0.98 ;
        RECT  0.54 0.82 0.70 2.22 ;
        RECT  0.54 1.94 0.90 2.22 ;
        RECT  2.26 0.68 2.42 2.14 ;
        RECT  0.54 2.06 1.50 2.22 ;
        RECT  1.34 2.06 1.50 2.54 ;
        RECT  2.14 1.86 2.30 2.54 ;
        RECT  1.34 2.38 2.30 2.54 ;
        RECT  3.10 0.68 3.46 0.96 ;
        RECT  3.10 0.68 3.26 2.14 ;
        RECT  3.10 1.86 3.46 2.14 ;
        RECT  4.22 0.68 4.62 0.96 ;
        RECT  4.46 1.16 4.82 1.44 ;
        RECT  4.46 0.68 4.62 2.14 ;
        RECT  4.22 1.86 4.62 2.14 ;
        RECT  2.66 0.68 2.94 0.96 ;
        RECT  4.78 0.72 5.14 1.00 ;
        RECT  2.72 0.68 2.88 2.14 ;
        RECT  2.66 1.86 2.94 2.14 ;
        RECT  4.98 0.72 5.14 2.20 ;
        RECT  4.78 1.92 5.14 2.20 ;
        RECT  2.78 1.86 2.94 2.46 ;
        RECT  4.78 1.92 4.94 2.46 ;
        RECT  2.78 2.30 4.94 2.46 ;
        RECT  5.86 0.72 6.16 1.00 ;
        RECT  5.86 0.72 6.02 2.20 ;
        RECT  5.82 1.92 6.10 2.20 ;
        RECT  5.30 0.72 5.58 1.00 ;
        RECT  6.66 1.48 6.94 1.76 ;
        RECT  6.26 1.60 6.94 1.76 ;
        RECT  5.36 0.72 5.52 2.20 ;
        RECT  5.30 1.92 5.58 2.20 ;
        RECT  5.42 1.92 5.58 2.52 ;
        RECT  6.26 1.60 6.42 2.52 ;
        RECT  5.42 2.36 6.42 2.52 ;
        RECT  6.92 0.72 7.26 1.00 ;
        RECT  6.18 1.16 7.26 1.32 ;
        RECT  6.18 1.16 6.46 1.44 ;
        RECT  7.10 0.72 7.26 2.20 ;
        RECT  7.10 1.92 7.38 2.20 ;
        RECT  7.60 0.44 9.08 0.60 ;
        RECT  8.80 0.44 9.08 0.80 ;
        RECT  7.48 0.76 7.76 1.04 ;
        RECT  7.60 0.44 7.76 2.20 ;
        RECT  7.60 1.92 7.90 2.20 ;
        RECT  8.62 0.96 8.90 1.24 ;
        RECT  8.62 1.46 9.56 1.62 ;
        RECT  9.28 1.40 9.56 1.68 ;
        RECT  8.62 0.96 8.78 2.12 ;
        RECT  8.62 1.84 8.90 2.12 ;
        RECT  8.00 0.76 8.30 1.04 ;
        RECT  9.66 0.96 9.94 1.24 ;
        RECT  9.66 1.84 9.94 2.12 ;
        RECT  8.14 0.76 8.30 2.20 ;
        RECT  8.26 1.92 8.42 2.44 ;
        RECT  9.75 0.96 9.91 2.70 ;
        RECT  8.26 2.28 9.91 2.44 ;
        RECT  9.75 2.42 10.04 2.70 ;
    END
END DFFDRBZSP2V1_0

MACRO DFFDRBZSP1V1_0
    CLASS CORE ;
    FOREIGN DFFDRBZSP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN TD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.62 1.86 3.94 2.14 ;
        RECT  3.62 1.42 3.78 2.14 ;
        RECT  3.42 1.42 3.78 1.70 ;
        END
    END TD
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.42 1.62 1.78 ;
        END
    END SEL
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 21.68  LAYER ME1  ;
        ANTENNADIFFAREA 9.16  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.60  LAYER ME1  ;
        ANTENNAMAXAREACAR 35.84  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.26 1.46 11.52 1.74 ;
        RECT  11.18 1.90 11.46 2.18 ;
        RECT  11.26 0.96 11.46 2.18 ;
        RECT  11.18 0.96 11.46 1.24 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 21.98  LAYER ME1  ;
        ANTENNADIFFAREA 9.16  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.60  LAYER ME1  ;
        ANTENNAMAXAREACAR 36.35  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.26 1.46 10.74 1.74 ;
        RECT  10.14 1.90 10.42 2.18 ;
        RECT  10.26 0.96 10.42 2.18 ;
        RECT  10.14 0.96 10.42 1.24 ;
        END
    END QB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.02 1.25 4.30 1.70 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END D
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.36 1.14 1.78 ;
        END
    END RB
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 11.60 0.28 ;
        RECT  11.14 -0.28 11.42 0.32 ;
        RECT  10.66 0.96 10.94 1.24 ;
        RECT  10.72 -0.28 10.88 1.24 ;
        RECT  9.14 0.96 9.42 1.24 ;
        RECT  9.24 -0.28 9.40 1.24 ;
        RECT  6.40 0.72 6.68 1.00 ;
        RECT  6.46 -0.28 6.62 1.00 ;
        RECT  3.70 0.68 3.98 0.96 ;
        RECT  3.76 -0.28 3.92 0.96 ;
        RECT  1.14 0.70 1.42 0.98 ;
        RECT  1.20 -0.28 1.36 0.98 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 11.60 3.48 ;
        RECT  11.14 2.88 11.42 3.48 ;
        RECT  10.66 1.90 10.94 2.18 ;
        RECT  10.72 1.90 10.88 3.48 ;
        RECT  9.14 2.62 9.42 3.48 ;
        RECT  6.58 1.92 6.86 2.20 ;
        RECT  6.64 1.92 6.80 3.48 ;
        RECT  3.70 2.62 3.98 3.48 ;
        RECT  0.92 2.62 1.20 3.48 ;
        RECT  0.10 1.94 0.38 2.22 ;
        RECT  0.16 1.94 0.32 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  1.66 0.70 1.94 0.98 ;
        RECT  1.78 1.20 2.10 1.48 ;
        RECT  1.78 0.70 1.94 2.22 ;
        RECT  1.66 1.94 1.94 2.22 ;
        RECT  0.10 0.70 0.38 0.98 ;
        RECT  2.14 0.68 2.42 0.96 ;
        RECT  0.10 0.82 0.70 0.98 ;
        RECT  0.54 0.82 0.70 2.22 ;
        RECT  0.54 1.94 0.90 2.22 ;
        RECT  2.26 0.68 2.42 2.14 ;
        RECT  0.54 2.06 1.50 2.22 ;
        RECT  1.34 2.06 1.50 2.54 ;
        RECT  2.14 1.86 2.30 2.54 ;
        RECT  1.34 2.38 2.30 2.54 ;
        RECT  3.10 0.68 3.46 0.96 ;
        RECT  3.10 0.68 3.26 2.14 ;
        RECT  3.10 1.86 3.46 2.14 ;
        RECT  4.22 0.68 4.62 0.96 ;
        RECT  4.46 1.16 4.82 1.44 ;
        RECT  4.46 0.68 4.62 2.14 ;
        RECT  4.22 1.86 4.62 2.14 ;
        RECT  2.66 0.68 2.94 0.96 ;
        RECT  4.78 0.72 5.14 1.00 ;
        RECT  2.72 0.68 2.88 2.14 ;
        RECT  2.66 1.86 2.94 2.14 ;
        RECT  4.98 0.72 5.14 2.20 ;
        RECT  4.78 1.92 5.14 2.20 ;
        RECT  2.78 1.86 2.94 2.46 ;
        RECT  4.78 1.92 4.94 2.46 ;
        RECT  2.78 2.30 4.94 2.46 ;
        RECT  5.86 0.72 6.16 1.00 ;
        RECT  5.86 0.72 6.02 2.20 ;
        RECT  5.82 1.92 6.10 2.20 ;
        RECT  5.30 0.72 5.58 1.00 ;
        RECT  6.66 1.48 6.94 1.76 ;
        RECT  6.26 1.60 6.94 1.76 ;
        RECT  5.36 0.72 5.52 2.20 ;
        RECT  5.30 1.92 5.58 2.20 ;
        RECT  5.42 1.92 5.58 2.52 ;
        RECT  6.26 1.60 6.42 2.52 ;
        RECT  5.42 2.36 6.42 2.52 ;
        RECT  6.92 0.72 7.26 1.00 ;
        RECT  6.18 1.16 7.26 1.32 ;
        RECT  6.18 1.16 6.46 1.44 ;
        RECT  7.10 0.72 7.26 2.20 ;
        RECT  7.10 1.92 7.38 2.20 ;
        RECT  7.60 0.44 9.08 0.60 ;
        RECT  8.80 0.44 9.08 0.80 ;
        RECT  7.48 0.76 7.76 1.04 ;
        RECT  7.60 0.44 7.76 2.20 ;
        RECT  7.60 1.92 7.90 2.20 ;
        RECT  8.62 0.96 8.90 1.24 ;
        RECT  8.62 1.46 9.56 1.62 ;
        RECT  9.28 1.40 9.56 1.68 ;
        RECT  8.62 0.96 8.78 2.12 ;
        RECT  8.62 1.84 8.90 2.12 ;
        RECT  8.00 0.76 8.30 1.04 ;
        RECT  9.66 0.96 9.94 1.24 ;
        RECT  9.66 1.84 9.94 2.12 ;
        RECT  8.14 0.76 8.30 2.20 ;
        RECT  8.26 1.92 8.42 2.44 ;
        RECT  9.75 0.96 9.91 2.70 ;
        RECT  8.26 2.28 9.91 2.44 ;
        RECT  9.75 2.42 10.04 2.70 ;
    END
END DFFDRBZSP1V1_0

MACRO DFFDRBSP8V1_1
    CLASS CORE ;
    FOREIGN DFFDRBSP8V1_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 22.68  LAYER ME1  ;
        ANTENNADIFFAREA 11.91  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.56  LAYER ME1  ;
        ANTENNAMAXAREACAR 14.59  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.32 1.84 11.60 2.12 ;
        RECT  11.32 0.96 11.60 1.24 ;
        RECT  11.32 0.96 11.48 2.12 ;
        RECT  10.40 1.52 11.48 1.68 ;
        RECT  10.40 1.46 10.74 1.74 ;
        RECT  10.28 1.84 10.56 2.12 ;
        RECT  10.40 0.96 10.56 2.12 ;
        RECT  10.28 0.96 10.56 1.24 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 22.68  LAYER ME1  ;
        ANTENNADIFFAREA 11.91  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.56  LAYER ME1  ;
        ANTENNAMAXAREACAR 14.59  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.24 1.84 9.52 2.12 ;
        RECT  9.24 0.96 9.52 1.24 ;
        RECT  9.24 0.96 9.40 2.12 ;
        RECT  8.06 1.52 9.40 1.68 ;
        RECT  8.20 1.84 8.48 2.12 ;
        RECT  8.20 0.96 8.48 1.24 ;
        RECT  8.20 0.96 8.36 2.12 ;
        RECT  8.06 1.46 8.36 1.74 ;
        END
    END Q
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.39 1.62 1.81 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END D
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.39 0.38 1.81 ;
        END
    END RB
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 12.40 0.28 ;
        RECT  11.90 -0.28 12.22 0.32 ;
        RECT  11.84 0.64 12.12 0.92 ;
        RECT  11.90 -0.28 12.06 0.92 ;
        RECT  10.80 0.64 11.08 0.92 ;
        RECT  10.86 -0.28 11.02 0.92 ;
        RECT  9.76 0.64 10.04 0.92 ;
        RECT  9.82 -0.28 9.98 0.92 ;
        RECT  8.72 0.64 9.00 0.92 ;
        RECT  8.78 -0.28 8.94 0.92 ;
        RECT  7.68 0.64 7.96 0.92 ;
        RECT  7.74 -0.28 7.90 0.92 ;
        RECT  6.68 0.96 6.96 1.24 ;
        RECT  6.78 -0.28 6.94 1.24 ;
        RECT  3.88 0.72 4.16 1.00 ;
        RECT  3.94 -0.28 4.10 1.00 ;
        RECT  1.14 0.68 1.42 0.96 ;
        RECT  1.20 -0.28 1.36 0.96 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 12.40 3.48 ;
        RECT  11.90 2.88 12.22 3.48 ;
        RECT  11.84 2.16 12.12 2.44 ;
        RECT  11.90 2.16 12.06 3.48 ;
        RECT  10.80 2.16 11.08 2.44 ;
        RECT  10.86 2.16 11.02 3.48 ;
        RECT  9.76 2.16 10.04 2.44 ;
        RECT  9.82 2.16 9.98 3.48 ;
        RECT  8.72 2.16 9.00 2.44 ;
        RECT  8.78 2.16 8.94 3.48 ;
        RECT  7.68 1.87 7.96 2.15 ;
        RECT  7.74 1.87 7.90 3.48 ;
        RECT  6.68 2.62 6.96 3.48 ;
        RECT  4.00 1.92 4.28 2.20 ;
        RECT  4.06 1.92 4.22 3.48 ;
        RECT  0.90 2.62 1.18 3.48 ;
        RECT  0.10 1.97 0.38 2.25 ;
        RECT  0.16 1.97 0.32 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  1.66 0.68 2.00 0.96 ;
        RECT  1.84 1.22 2.16 1.50 ;
        RECT  1.84 0.68 2.00 2.25 ;
        RECT  1.66 1.97 2.00 2.25 ;
        RECT  0.10 0.68 0.38 0.96 ;
        RECT  0.10 0.80 0.70 0.96 ;
        RECT  2.20 0.72 2.48 1.00 ;
        RECT  0.54 0.80 0.70 2.25 ;
        RECT  0.54 1.97 0.90 2.25 ;
        RECT  2.32 0.72 2.48 2.20 ;
        RECT  0.54 2.09 1.50 2.25 ;
        RECT  1.34 2.09 1.50 2.57 ;
        RECT  2.20 1.92 2.36 2.57 ;
        RECT  1.34 2.41 2.36 2.57 ;
        RECT  3.28 0.72 3.59 1.00 ;
        RECT  3.28 0.72 3.44 2.20 ;
        RECT  3.24 1.92 3.52 2.20 ;
        RECT  2.72 0.72 3.00 1.00 ;
        RECT  4.08 1.48 4.36 1.76 ;
        RECT  3.68 1.60 4.36 1.76 ;
        RECT  2.78 0.72 2.94 2.20 ;
        RECT  2.72 1.92 3.00 2.20 ;
        RECT  2.84 1.92 3.00 2.52 ;
        RECT  3.68 1.60 3.84 2.52 ;
        RECT  2.84 2.36 3.84 2.52 ;
        RECT  4.40 0.72 4.68 1.00 ;
        RECT  3.60 1.16 4.68 1.32 ;
        RECT  3.60 1.16 3.88 1.44 ;
        RECT  4.52 0.72 4.68 2.20 ;
        RECT  4.52 1.92 4.80 2.20 ;
        RECT  5.16 0.44 6.62 0.60 ;
        RECT  6.34 0.44 6.62 0.80 ;
        RECT  5.16 0.44 5.32 1.04 ;
        RECT  5.04 0.76 5.32 1.04 ;
        RECT  5.10 0.76 5.26 2.20 ;
        RECT  5.04 1.92 5.32 2.20 ;
        RECT  6.16 0.96 6.44 1.24 ;
        RECT  6.16 1.46 7.16 1.62 ;
        RECT  6.88 1.40 7.16 1.68 ;
        RECT  6.16 0.96 6.32 2.12 ;
        RECT  6.16 1.84 6.44 2.12 ;
        RECT  5.56 0.76 5.84 1.04 ;
        RECT  7.20 0.96 7.48 1.24 ;
        RECT  7.20 1.84 7.48 2.12 ;
        RECT  5.62 0.76 5.78 2.20 ;
        RECT  5.56 1.92 5.84 2.20 ;
        RECT  5.68 1.92 5.84 2.44 ;
        RECT  7.32 0.96 7.48 2.70 ;
        RECT  5.68 2.28 7.48 2.44 ;
        RECT  7.30 2.42 7.58 2.70 ;
    END
END DFFDRBSP8V1_1

MACRO DFFDRBSP8V1_0
    CLASS CORE ;
    FOREIGN DFFDRBSP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.30 1.12 2.72 1.40 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.46 1.39 0.74 1.81 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 23.36  LAYER ME1  ;
        ANTENNADIFFAREA 12.07  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.79  LAYER ME1  ;
        ANTENNAMAXAREACAR 13.05  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.64 1.84 9.92 2.12 ;
        RECT  9.64 0.96 9.92 1.24 ;
        RECT  9.64 0.96 9.80 2.12 ;
        RECT  8.46 1.52 9.80 1.68 ;
        RECT  8.60 1.84 8.88 2.12 ;
        RECT  8.60 0.96 8.88 1.24 ;
        RECT  8.60 0.96 8.76 2.12 ;
        RECT  8.46 1.46 8.76 1.74 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 23.36  LAYER ME1  ;
        ANTENNADIFFAREA 11.87  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.79  LAYER ME1  ;
        ANTENNAMAXAREACAR 13.05  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.72 1.84 12.00 2.12 ;
        RECT  11.72 0.96 12.00 1.24 ;
        RECT  11.72 0.96 11.88 2.12 ;
        RECT  10.80 1.52 11.88 1.68 ;
        RECT  10.68 1.84 10.96 2.12 ;
        RECT  10.80 0.96 10.96 2.12 ;
        RECT  10.68 0.96 10.96 1.24 ;
        END
    END QB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.64 1.12 2.06 1.40 ;
        END
    END RB
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 12.80 0.28 ;
        RECT  12.30 -0.28 12.62 0.32 ;
        RECT  12.24 0.64 12.52 0.92 ;
        RECT  12.30 -0.28 12.46 0.92 ;
        RECT  11.20 0.64 11.48 0.92 ;
        RECT  11.26 -0.28 11.42 0.92 ;
        RECT  10.16 0.64 10.44 0.92 ;
        RECT  10.22 -0.28 10.38 0.92 ;
        RECT  9.12 0.64 9.40 0.92 ;
        RECT  9.18 -0.28 9.34 0.92 ;
        RECT  8.08 0.64 8.36 0.92 ;
        RECT  8.14 -0.28 8.30 0.92 ;
        RECT  7.08 0.96 7.36 1.24 ;
        RECT  7.18 -0.28 7.34 1.24 ;
        RECT  4.36 0.68 4.64 0.96 ;
        RECT  4.42 -0.28 4.58 0.96 ;
        RECT  1.64 0.68 1.92 0.96 ;
        RECT  1.70 -0.28 1.86 0.96 ;
        RECT  0.62 0.50 0.90 0.78 ;
        RECT  0.68 -0.28 0.84 0.78 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 12.80 3.48 ;
        RECT  12.30 2.88 12.62 3.48 ;
        RECT  12.24 2.16 12.52 2.44 ;
        RECT  12.30 2.16 12.46 3.48 ;
        RECT  11.20 2.16 11.48 2.44 ;
        RECT  11.26 2.16 11.42 3.48 ;
        RECT  10.16 2.16 10.44 2.44 ;
        RECT  10.22 2.16 10.38 3.48 ;
        RECT  9.12 2.16 9.40 2.44 ;
        RECT  9.18 2.16 9.34 3.48 ;
        RECT  8.08 1.87 8.36 2.15 ;
        RECT  8.14 1.87 8.30 3.48 ;
        RECT  7.08 2.62 7.36 3.48 ;
        RECT  4.52 1.92 4.80 2.20 ;
        RECT  4.58 1.92 4.74 3.48 ;
        RECT  2.16 1.92 2.44 2.20 ;
        RECT  2.24 1.92 2.40 3.48 ;
        RECT  0.62 1.97 0.90 2.25 ;
        RECT  0.68 1.97 0.84 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.08 0.50 0.38 0.78 ;
        RECT  0.08 1.00 1.16 1.16 ;
        RECT  0.88 0.94 1.16 1.22 ;
        RECT  0.08 0.50 0.24 2.25 ;
        RECT  0.08 1.97 0.38 2.25 ;
        RECT  1.14 0.50 1.48 0.78 ;
        RECT  1.14 1.97 1.48 2.25 ;
        RECT  1.32 0.50 1.48 2.70 ;
        RECT  1.28 2.42 1.56 2.70 ;
        RECT  2.68 0.68 3.04 0.96 ;
        RECT  1.76 1.60 3.04 1.76 ;
        RECT  1.76 1.60 1.92 2.20 ;
        RECT  1.64 1.92 1.92 2.20 ;
        RECT  2.88 0.68 3.04 2.20 ;
        RECT  2.68 1.92 3.04 2.20 ;
        RECT  3.20 0.68 3.48 0.96 ;
        RECT  3.26 0.68 3.42 2.20 ;
        RECT  3.20 1.92 3.48 2.20 ;
        RECT  3.32 1.92 3.48 2.70 ;
        RECT  3.86 2.42 4.14 2.70 ;
        RECT  3.32 2.54 4.14 2.70 ;
        RECT  3.72 0.68 4.08 0.96 ;
        RECT  3.92 0.68 4.08 2.20 ;
        RECT  3.86 1.92 4.14 2.20 ;
        RECT  4.88 0.68 5.20 0.96 ;
        RECT  4.38 1.44 5.20 1.60 ;
        RECT  4.38 1.38 4.66 1.66 ;
        RECT  5.04 0.68 5.20 2.20 ;
        RECT  5.04 1.92 5.32 2.20 ;
        RECT  5.56 0.44 7.02 0.60 ;
        RECT  6.74 0.44 7.02 0.80 ;
        RECT  5.44 0.76 5.72 1.04 ;
        RECT  5.56 0.44 5.72 2.20 ;
        RECT  5.56 1.92 5.84 2.20 ;
        RECT  6.56 0.96 6.84 1.24 ;
        RECT  6.56 1.46 7.56 1.62 ;
        RECT  7.28 1.40 7.56 1.68 ;
        RECT  6.56 0.96 6.72 2.12 ;
        RECT  6.56 1.84 6.84 2.12 ;
        RECT  5.96 0.76 6.24 1.04 ;
        RECT  7.60 0.96 7.88 1.24 ;
        RECT  7.60 1.84 7.88 2.12 ;
        RECT  6.08 0.76 6.24 2.20 ;
        RECT  6.20 1.92 6.36 2.44 ;
        RECT  7.72 0.96 7.88 2.70 ;
        RECT  6.20 2.28 7.88 2.44 ;
        RECT  7.70 2.42 7.98 2.70 ;
    END
END DFFDRBSP8V1_0

MACRO DFFDRBSP4V1_1
    CLASS CORE ;
    FOREIGN DFFDRBSP4V1_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.39 0.38 1.81 ;
        END
    END RB
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.39 1.62 1.81 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 19.14  LAYER ME1  ;
        ANTENNADIFFAREA 9.14  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.98  LAYER ME1  ;
        ANTENNAMAXAREACAR 19.55  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.26 1.46 9.54 1.74 ;
        RECT  9.24 1.84 9.52 2.12 ;
        RECT  9.26 0.96 9.52 2.12 ;
        RECT  9.24 0.96 9.52 1.24 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 18.85  LAYER ME1  ;
        ANTENNADIFFAREA 9.14  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.98  LAYER ME1  ;
        ANTENNAMAXAREACAR 19.25  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.20 1.84 8.48 2.12 ;
        RECT  8.20 0.96 8.48 1.24 ;
        RECT  8.20 0.96 8.36 2.12 ;
        RECT  8.06 1.46 8.36 1.74 ;
        END
    END Q
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 10.40 3.48 ;
        RECT  9.82 2.88 10.22 3.48 ;
        RECT  9.76 2.16 10.04 2.44 ;
        RECT  9.82 2.16 9.98 3.48 ;
        RECT  8.72 2.16 9.00 2.44 ;
        RECT  8.78 2.16 8.94 3.48 ;
        RECT  7.68 1.87 7.96 2.15 ;
        RECT  7.74 1.87 7.90 3.48 ;
        RECT  6.68 2.62 6.96 3.48 ;
        RECT  4.00 1.92 4.28 2.20 ;
        RECT  4.06 1.92 4.22 3.48 ;
        RECT  0.90 2.62 1.18 3.48 ;
        RECT  0.10 1.97 0.38 2.25 ;
        RECT  0.16 1.97 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 10.40 0.28 ;
        RECT  9.82 -0.28 10.22 0.32 ;
        RECT  9.76 0.64 10.04 0.92 ;
        RECT  9.82 -0.28 9.98 0.92 ;
        RECT  8.72 0.64 9.00 0.92 ;
        RECT  8.78 -0.28 8.94 0.92 ;
        RECT  7.68 0.64 7.96 0.92 ;
        RECT  7.74 -0.28 7.90 0.92 ;
        RECT  6.68 0.96 6.96 1.24 ;
        RECT  6.78 -0.28 6.94 1.24 ;
        RECT  3.88 0.72 4.16 1.00 ;
        RECT  3.94 -0.28 4.10 1.00 ;
        RECT  1.14 0.68 1.42 0.96 ;
        RECT  1.20 -0.28 1.36 0.96 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  1.66 0.68 2.00 0.96 ;
        RECT  1.84 1.22 2.16 1.50 ;
        RECT  1.84 0.68 2.00 2.25 ;
        RECT  1.66 1.97 2.00 2.25 ;
        RECT  0.10 0.68 0.38 0.96 ;
        RECT  0.10 0.80 0.70 0.96 ;
        RECT  2.20 0.72 2.48 1.00 ;
        RECT  0.54 0.80 0.70 2.25 ;
        RECT  0.54 1.97 0.90 2.25 ;
        RECT  2.32 0.72 2.48 2.20 ;
        RECT  0.54 2.09 1.50 2.25 ;
        RECT  1.34 2.09 1.50 2.57 ;
        RECT  2.20 1.92 2.36 2.57 ;
        RECT  1.34 2.41 2.36 2.57 ;
        RECT  3.28 0.72 3.59 1.00 ;
        RECT  3.28 0.72 3.44 2.20 ;
        RECT  3.24 1.92 3.52 2.20 ;
        RECT  2.72 0.72 3.00 1.00 ;
        RECT  4.08 1.48 4.36 1.76 ;
        RECT  3.68 1.60 4.36 1.76 ;
        RECT  2.78 0.72 2.94 2.20 ;
        RECT  2.72 1.92 3.00 2.20 ;
        RECT  2.84 1.92 3.00 2.52 ;
        RECT  3.68 1.60 3.84 2.52 ;
        RECT  2.84 2.36 3.84 2.52 ;
        RECT  4.40 0.72 4.68 1.00 ;
        RECT  3.60 1.16 4.68 1.32 ;
        RECT  3.60 1.16 3.88 1.44 ;
        RECT  4.52 0.72 4.68 2.20 ;
        RECT  4.52 1.92 4.80 2.20 ;
        RECT  5.16 0.44 6.62 0.60 ;
        RECT  6.34 0.44 6.62 0.80 ;
        RECT  5.16 0.44 5.32 1.04 ;
        RECT  5.04 0.76 5.32 1.04 ;
        RECT  5.10 0.76 5.26 2.20 ;
        RECT  5.04 1.92 5.32 2.20 ;
        RECT  6.16 0.96 6.44 1.24 ;
        RECT  6.16 1.46 7.16 1.62 ;
        RECT  6.88 1.40 7.16 1.68 ;
        RECT  6.16 0.96 6.32 2.12 ;
        RECT  6.16 1.84 6.44 2.12 ;
        RECT  5.56 0.76 5.84 1.04 ;
        RECT  7.20 0.96 7.48 1.24 ;
        RECT  7.20 1.84 7.48 2.12 ;
        RECT  5.62 0.76 5.78 2.20 ;
        RECT  5.56 1.92 5.84 2.20 ;
        RECT  5.68 1.92 5.84 2.44 ;
        RECT  7.32 0.96 7.48 2.70 ;
        RECT  5.68 2.28 7.48 2.44 ;
        RECT  7.30 2.42 7.58 2.70 ;
    END
END DFFDRBSP4V1_1

MACRO DFFDRBSP4V1_0
    CLASS CORE ;
    FOREIGN DFFDRBSP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.64 1.12 2.06 1.40 ;
        END
    END RB
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 19.52  LAYER ME1  ;
        ANTENNADIFFAREA 9.31  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.21  LAYER ME1  ;
        ANTENNAMAXAREACAR 16.08  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.64 1.84 9.92 2.12 ;
        RECT  9.64 0.96 9.92 1.24 ;
        RECT  9.72 0.96 9.88 2.12 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 19.78  LAYER ME1  ;
        ANTENNADIFFAREA 9.31  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.21  LAYER ME1  ;
        ANTENNAMAXAREACAR 16.28  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.60 1.84 8.88 2.12 ;
        RECT  8.60 0.96 8.88 1.24 ;
        RECT  8.60 0.96 8.76 2.12 ;
        RECT  8.46 1.46 8.76 1.74 ;
        END
    END Q
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.46 1.39 0.74 1.81 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.30 1.12 2.72 1.40 ;
        END
    END D
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 10.80 3.48 ;
        RECT  10.22 2.88 10.62 3.48 ;
        RECT  10.16 2.16 10.44 2.44 ;
        RECT  10.22 2.16 10.38 3.48 ;
        RECT  9.12 2.16 9.40 2.44 ;
        RECT  9.18 2.16 9.34 3.48 ;
        RECT  8.08 1.87 8.36 2.15 ;
        RECT  8.14 1.87 8.30 3.48 ;
        RECT  7.08 2.62 7.36 3.48 ;
        RECT  4.52 1.92 4.80 2.20 ;
        RECT  4.58 1.92 4.74 3.48 ;
        RECT  2.16 1.92 2.44 2.20 ;
        RECT  2.24 1.92 2.40 3.48 ;
        RECT  0.62 1.97 0.90 2.25 ;
        RECT  0.68 1.97 0.84 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 10.80 0.28 ;
        RECT  10.22 -0.28 10.62 0.32 ;
        RECT  10.16 0.64 10.44 0.92 ;
        RECT  10.22 -0.28 10.38 0.92 ;
        RECT  9.12 0.64 9.40 0.92 ;
        RECT  9.18 -0.28 9.34 0.92 ;
        RECT  8.08 0.64 8.36 0.92 ;
        RECT  8.14 -0.28 8.30 0.92 ;
        RECT  7.08 0.96 7.36 1.24 ;
        RECT  7.18 -0.28 7.34 1.24 ;
        RECT  4.36 0.68 4.64 0.96 ;
        RECT  4.42 -0.28 4.58 0.96 ;
        RECT  1.64 0.68 1.92 0.96 ;
        RECT  1.70 -0.28 1.86 0.96 ;
        RECT  0.62 0.50 0.90 0.78 ;
        RECT  0.68 -0.28 0.84 0.78 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.08 0.50 0.38 0.78 ;
        RECT  0.08 1.00 1.16 1.16 ;
        RECT  0.88 0.94 1.16 1.22 ;
        RECT  0.08 0.50 0.24 2.25 ;
        RECT  0.08 1.97 0.38 2.25 ;
        RECT  1.14 0.50 1.48 0.78 ;
        RECT  1.14 1.97 1.48 2.25 ;
        RECT  1.32 0.50 1.48 2.70 ;
        RECT  1.28 2.42 1.56 2.70 ;
        RECT  2.68 0.68 3.04 0.96 ;
        RECT  1.76 1.60 3.04 1.76 ;
        RECT  1.76 1.60 1.92 2.20 ;
        RECT  1.64 1.92 1.92 2.20 ;
        RECT  2.88 0.68 3.04 2.20 ;
        RECT  2.68 1.92 3.04 2.20 ;
        RECT  3.20 0.68 3.48 0.96 ;
        RECT  3.26 0.68 3.42 2.20 ;
        RECT  3.20 1.92 3.48 2.20 ;
        RECT  3.32 1.92 3.48 2.70 ;
        RECT  3.86 2.42 4.14 2.70 ;
        RECT  3.32 2.54 4.14 2.70 ;
        RECT  3.72 0.68 4.08 0.96 ;
        RECT  3.92 0.68 4.08 2.20 ;
        RECT  3.86 1.92 4.14 2.20 ;
        RECT  4.88 0.68 5.20 0.96 ;
        RECT  4.38 1.44 5.20 1.60 ;
        RECT  4.38 1.38 4.66 1.66 ;
        RECT  5.04 0.68 5.20 2.20 ;
        RECT  5.04 1.92 5.32 2.20 ;
        RECT  5.56 0.44 7.02 0.60 ;
        RECT  6.74 0.44 7.02 0.80 ;
        RECT  5.44 0.76 5.72 1.04 ;
        RECT  5.56 0.44 5.72 2.20 ;
        RECT  5.56 1.92 5.84 2.20 ;
        RECT  6.56 0.96 6.84 1.24 ;
        RECT  6.56 1.46 7.56 1.62 ;
        RECT  7.28 1.40 7.56 1.68 ;
        RECT  6.56 0.96 6.72 2.12 ;
        RECT  6.56 1.84 6.84 2.12 ;
        RECT  5.96 0.76 6.24 1.04 ;
        RECT  7.60 0.96 7.88 1.24 ;
        RECT  7.60 1.84 7.88 2.12 ;
        RECT  6.08 0.76 6.24 2.20 ;
        RECT  6.20 1.92 6.36 2.44 ;
        RECT  7.72 0.96 7.88 2.70 ;
        RECT  6.20 2.28 7.88 2.44 ;
        RECT  7.70 2.42 7.98 2.70 ;
    END
END DFFDRBSP4V1_0

MACRO DFFDRBSP2V1_1
    CLASS CORE ;
    FOREIGN DFFDRBSP2V1_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 17.17  LAYER ME1  ;
        ANTENNADIFFAREA 7.80  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.69  LAYER ME1  ;
        ANTENNAMAXAREACAR 24.84  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.68 1.84 7.96 2.12 ;
        RECT  7.68 0.96 7.96 1.24 ;
        RECT  7.68 0.96 7.94 2.12 ;
        RECT  7.66 1.46 7.94 1.74 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 16.88  LAYER ME1  ;
        ANTENNADIFFAREA 7.80  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.69  LAYER ME1  ;
        ANTENNAMAXAREACAR 24.43  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.84 1.46 9.12 1.74 ;
        RECT  8.72 1.84 9.00 2.12 ;
        RECT  8.84 0.96 9.00 2.12 ;
        RECT  8.72 0.96 9.00 1.24 ;
        END
    END QB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.39 1.62 1.81 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END D
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.39 0.38 1.81 ;
        END
    END RB
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 9.20 0.28 ;
        RECT  8.74 -0.28 9.02 0.32 ;
        RECT  8.20 0.64 8.48 0.92 ;
        RECT  8.26 -0.28 8.42 0.92 ;
        RECT  6.68 0.96 6.96 1.24 ;
        RECT  6.78 -0.28 6.94 1.24 ;
        RECT  3.88 0.72 4.16 1.00 ;
        RECT  3.94 -0.28 4.10 1.00 ;
        RECT  1.14 0.68 1.42 0.96 ;
        RECT  1.20 -0.28 1.36 0.96 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 9.20 3.48 ;
        RECT  8.74 2.88 9.02 3.48 ;
        RECT  8.20 2.16 8.48 2.44 ;
        RECT  8.26 2.16 8.42 3.48 ;
        RECT  6.68 2.62 6.96 3.48 ;
        RECT  4.00 1.92 4.28 2.20 ;
        RECT  4.06 1.92 4.22 3.48 ;
        RECT  0.90 2.62 1.18 3.48 ;
        RECT  0.10 1.97 0.38 2.25 ;
        RECT  0.16 1.97 0.32 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  1.66 0.68 2.00 0.96 ;
        RECT  1.84 1.22 2.16 1.50 ;
        RECT  1.84 0.68 2.00 2.25 ;
        RECT  1.66 1.97 2.00 2.25 ;
        RECT  0.10 0.68 0.38 0.96 ;
        RECT  0.10 0.80 0.70 0.96 ;
        RECT  2.20 0.72 2.48 1.00 ;
        RECT  0.54 0.80 0.70 2.25 ;
        RECT  0.54 1.97 0.90 2.25 ;
        RECT  2.32 0.72 2.48 2.20 ;
        RECT  0.54 2.09 1.50 2.25 ;
        RECT  1.34 2.09 1.50 2.57 ;
        RECT  2.20 1.92 2.36 2.57 ;
        RECT  1.34 2.41 2.36 2.57 ;
        RECT  3.28 0.72 3.59 1.00 ;
        RECT  3.28 0.72 3.44 2.20 ;
        RECT  3.24 1.92 3.52 2.20 ;
        RECT  2.72 0.72 3.00 1.00 ;
        RECT  4.08 1.48 4.36 1.76 ;
        RECT  3.68 1.60 4.36 1.76 ;
        RECT  2.78 0.72 2.94 2.20 ;
        RECT  2.72 1.92 3.00 2.20 ;
        RECT  2.84 1.92 3.00 2.52 ;
        RECT  3.68 1.60 3.84 2.52 ;
        RECT  2.84 2.36 3.84 2.52 ;
        RECT  4.40 0.72 4.68 1.00 ;
        RECT  3.60 1.16 4.68 1.32 ;
        RECT  3.60 1.16 3.88 1.44 ;
        RECT  4.52 0.72 4.68 2.20 ;
        RECT  4.52 1.92 4.80 2.20 ;
        RECT  5.16 0.44 6.62 0.60 ;
        RECT  6.34 0.44 6.62 0.80 ;
        RECT  5.16 0.44 5.32 1.04 ;
        RECT  5.04 0.76 5.32 1.04 ;
        RECT  5.10 0.76 5.26 2.20 ;
        RECT  5.04 1.92 5.32 2.20 ;
        RECT  6.16 0.96 6.44 1.24 ;
        RECT  6.16 1.46 7.16 1.62 ;
        RECT  6.88 1.40 7.16 1.68 ;
        RECT  6.16 0.96 6.32 2.12 ;
        RECT  6.16 1.84 6.44 2.12 ;
        RECT  5.56 0.76 5.84 1.04 ;
        RECT  7.20 0.96 7.48 1.24 ;
        RECT  7.20 1.84 7.48 2.12 ;
        RECT  5.62 0.76 5.78 2.20 ;
        RECT  5.56 1.92 5.84 2.20 ;
        RECT  5.68 1.92 5.84 2.44 ;
        RECT  7.32 0.96 7.48 2.70 ;
        RECT  5.68 2.28 7.48 2.44 ;
        RECT  7.30 2.42 7.58 2.70 ;
    END
END DFFDRBSP2V1_1

MACRO DFFDRBSP2V1_0
    CLASS CORE ;
    FOREIGN DFFDRBSP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.30 1.12 2.72 1.40 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.46 1.39 0.74 1.81 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 17.56  LAYER ME1  ;
        ANTENNADIFFAREA 7.96  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.93  LAYER ME1  ;
        ANTENNAMAXAREACAR 18.95  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.08 1.84 8.36 2.12 ;
        RECT  8.08 0.96 8.36 1.24 ;
        RECT  8.12 0.96 8.28 2.12 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 17.81  LAYER ME1  ;
        ANTENNADIFFAREA 7.96  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.93  LAYER ME1  ;
        ANTENNAMAXAREACAR 19.23  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.12 1.84 9.48 2.12 ;
        RECT  9.32 0.96 9.48 2.12 ;
        RECT  9.12 0.96 9.48 1.24 ;
        END
    END QB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.64 1.12 2.06 1.40 ;
        END
    END RB
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 9.60 0.28 ;
        RECT  9.14 -0.28 9.42 0.32 ;
        RECT  8.60 0.64 8.88 0.92 ;
        RECT  8.66 -0.28 8.82 0.92 ;
        RECT  7.08 0.96 7.36 1.24 ;
        RECT  7.18 -0.28 7.34 1.24 ;
        RECT  4.36 0.68 4.64 0.96 ;
        RECT  4.42 -0.28 4.58 0.96 ;
        RECT  1.64 0.68 1.92 0.96 ;
        RECT  1.70 -0.28 1.86 0.96 ;
        RECT  0.62 0.50 0.90 0.78 ;
        RECT  0.68 -0.28 0.84 0.78 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 9.60 3.48 ;
        RECT  9.14 2.88 9.42 3.48 ;
        RECT  8.60 2.16 8.88 2.44 ;
        RECT  8.66 2.16 8.82 3.48 ;
        RECT  7.08 2.62 7.36 3.48 ;
        RECT  4.52 1.92 4.80 2.20 ;
        RECT  4.58 1.92 4.74 3.48 ;
        RECT  2.16 1.92 2.44 2.20 ;
        RECT  2.24 1.92 2.40 3.48 ;
        RECT  0.62 1.97 0.90 2.25 ;
        RECT  0.68 1.97 0.84 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.08 0.50 0.38 0.78 ;
        RECT  0.08 1.00 1.16 1.16 ;
        RECT  0.88 0.94 1.16 1.22 ;
        RECT  0.08 0.50 0.24 2.25 ;
        RECT  0.08 1.97 0.38 2.25 ;
        RECT  1.14 0.50 1.48 0.78 ;
        RECT  1.14 1.97 1.48 2.25 ;
        RECT  1.32 0.50 1.48 2.70 ;
        RECT  1.28 2.42 1.56 2.70 ;
        RECT  2.68 0.68 3.04 0.96 ;
        RECT  1.76 1.60 3.04 1.76 ;
        RECT  1.76 1.60 1.92 2.20 ;
        RECT  1.64 1.92 1.92 2.20 ;
        RECT  2.88 0.68 3.04 2.20 ;
        RECT  2.68 1.92 3.04 2.20 ;
        RECT  3.20 0.68 3.48 0.96 ;
        RECT  3.26 0.68 3.42 2.20 ;
        RECT  3.20 1.92 3.48 2.20 ;
        RECT  3.32 1.92 3.48 2.70 ;
        RECT  3.86 2.42 4.14 2.70 ;
        RECT  3.32 2.54 4.14 2.70 ;
        RECT  3.72 0.68 4.08 0.96 ;
        RECT  3.92 0.68 4.08 2.20 ;
        RECT  3.86 1.92 4.14 2.20 ;
        RECT  4.88 0.68 5.20 0.96 ;
        RECT  4.38 1.44 5.20 1.60 ;
        RECT  4.38 1.38 4.66 1.66 ;
        RECT  5.04 0.68 5.20 2.20 ;
        RECT  5.04 1.92 5.32 2.20 ;
        RECT  5.56 0.44 7.02 0.60 ;
        RECT  6.74 0.44 7.02 0.80 ;
        RECT  5.44 0.76 5.72 1.04 ;
        RECT  5.56 0.44 5.72 2.20 ;
        RECT  5.56 1.92 5.84 2.20 ;
        RECT  6.56 0.96 6.84 1.24 ;
        RECT  6.56 1.46 7.56 1.62 ;
        RECT  7.28 1.40 7.56 1.68 ;
        RECT  6.56 0.96 6.72 2.12 ;
        RECT  6.56 1.84 6.84 2.12 ;
        RECT  5.96 0.76 6.24 1.04 ;
        RECT  7.60 0.96 7.88 1.24 ;
        RECT  7.60 1.84 7.88 2.12 ;
        RECT  6.08 0.76 6.24 2.20 ;
        RECT  6.20 1.92 6.36 2.44 ;
        RECT  7.72 0.96 7.88 2.70 ;
        RECT  6.20 2.28 7.88 2.44 ;
        RECT  7.70 2.42 7.98 2.70 ;
    END
END DFFDRBSP2V1_0

MACRO DFFDRBSP1V1_1
    CLASS CORE ;
    FOREIGN DFFDRBSP1V1_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.39 1.62 1.81 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 16.98  LAYER ME1  ;
        ANTENNADIFFAREA 7.11  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.54  LAYER ME1  ;
        ANTENNAMAXAREACAR 31.59  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.84 1.46 9.12 1.74 ;
        RECT  8.72 1.84 9.00 2.12 ;
        RECT  8.84 0.96 9.00 2.12 ;
        RECT  8.72 0.96 9.00 1.24 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 17.27  LAYER ME1  ;
        ANTENNADIFFAREA 7.11  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.54  LAYER ME1  ;
        ANTENNAMAXAREACAR 32.12  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.68 1.84 7.96 2.12 ;
        RECT  7.68 0.96 7.96 1.24 ;
        RECT  7.68 0.96 7.94 2.12 ;
        RECT  7.66 1.46 7.94 1.74 ;
        END
    END Q
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.39 0.38 1.81 ;
        END
    END RB
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 9.20 3.48 ;
        RECT  8.74 2.88 9.02 3.48 ;
        RECT  8.20 1.84 8.48 2.12 ;
        RECT  8.26 1.84 8.42 3.48 ;
        RECT  6.68 2.62 6.96 3.48 ;
        RECT  4.00 1.92 4.28 2.20 ;
        RECT  4.06 1.92 4.22 3.48 ;
        RECT  0.90 2.62 1.18 3.48 ;
        RECT  0.10 1.97 0.38 2.25 ;
        RECT  0.16 1.97 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 9.20 0.28 ;
        RECT  8.74 -0.28 9.02 0.32 ;
        RECT  8.20 0.96 8.48 1.24 ;
        RECT  8.26 -0.28 8.42 1.24 ;
        RECT  6.68 0.96 6.96 1.24 ;
        RECT  6.78 -0.28 6.94 1.24 ;
        RECT  3.88 0.72 4.16 1.00 ;
        RECT  3.94 -0.28 4.10 1.00 ;
        RECT  1.14 0.68 1.42 0.96 ;
        RECT  1.20 -0.28 1.36 0.96 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  1.66 0.68 2.00 0.96 ;
        RECT  1.84 1.22 2.16 1.50 ;
        RECT  1.84 0.68 2.00 2.25 ;
        RECT  1.66 1.97 2.00 2.25 ;
        RECT  0.10 0.68 0.38 0.96 ;
        RECT  0.10 0.80 0.70 0.96 ;
        RECT  2.20 0.72 2.48 1.00 ;
        RECT  0.54 0.80 0.70 2.25 ;
        RECT  0.54 1.97 0.90 2.25 ;
        RECT  2.32 0.72 2.48 2.20 ;
        RECT  0.54 2.09 1.50 2.25 ;
        RECT  1.34 2.09 1.50 2.57 ;
        RECT  2.20 1.92 2.36 2.57 ;
        RECT  1.34 2.41 2.36 2.57 ;
        RECT  3.28 0.72 3.59 1.00 ;
        RECT  3.28 0.72 3.44 2.20 ;
        RECT  3.24 1.92 3.52 2.20 ;
        RECT  2.72 0.72 3.00 1.00 ;
        RECT  4.08 1.48 4.36 1.76 ;
        RECT  3.68 1.60 4.36 1.76 ;
        RECT  2.78 0.72 2.94 2.20 ;
        RECT  2.72 1.92 3.00 2.20 ;
        RECT  2.84 1.92 3.00 2.52 ;
        RECT  3.68 1.60 3.84 2.52 ;
        RECT  2.84 2.36 3.84 2.52 ;
        RECT  4.40 0.72 4.68 1.00 ;
        RECT  3.60 1.16 4.68 1.32 ;
        RECT  3.60 1.16 3.88 1.44 ;
        RECT  4.52 0.72 4.68 2.20 ;
        RECT  4.52 1.92 4.80 2.20 ;
        RECT  5.16 0.44 6.62 0.60 ;
        RECT  6.34 0.44 6.62 0.80 ;
        RECT  5.16 0.44 5.32 1.04 ;
        RECT  5.04 0.76 5.32 1.04 ;
        RECT  5.10 0.76 5.26 2.20 ;
        RECT  5.04 1.92 5.32 2.20 ;
        RECT  6.16 0.96 6.44 1.24 ;
        RECT  6.16 1.46 7.16 1.62 ;
        RECT  6.88 1.40 7.16 1.68 ;
        RECT  6.16 0.96 6.32 2.12 ;
        RECT  6.16 1.84 6.44 2.12 ;
        RECT  5.56 0.76 5.84 1.04 ;
        RECT  7.20 0.96 7.48 1.24 ;
        RECT  7.20 1.84 7.48 2.12 ;
        RECT  5.62 0.76 5.78 2.20 ;
        RECT  5.56 1.92 5.84 2.20 ;
        RECT  5.68 1.92 5.84 2.44 ;
        RECT  7.32 0.96 7.48 2.44 ;
        RECT  5.68 2.28 7.62 2.44 ;
        RECT  7.34 2.28 7.62 2.62 ;
    END
END DFFDRBSP1V1_1

MACRO DFFDRBSP1V1_0
    CLASS CORE ;
    FOREIGN DFFDRBSP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 17.93  LAYER ME1  ;
        ANTENNADIFFAREA 7.27  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.77  LAYER ME1  ;
        ANTENNAMAXAREACAR 23.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.12 1.84 9.48 2.12 ;
        RECT  9.32 0.96 9.48 2.12 ;
        RECT  9.12 0.96 9.48 1.24 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 17.68  LAYER ME1  ;
        ANTENNADIFFAREA 7.27  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.77  LAYER ME1  ;
        ANTENNAMAXAREACAR 22.87  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.08 1.84 8.36 2.12 ;
        RECT  8.08 0.96 8.36 1.24 ;
        RECT  8.12 0.96 8.28 2.12 ;
        END
    END Q
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.46 1.39 0.74 1.81 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.30 1.12 2.72 1.40 ;
        END
    END D
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.64 1.12 2.06 1.40 ;
        END
    END RB
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 9.60 3.48 ;
        RECT  9.14 2.88 9.42 3.48 ;
        RECT  8.60 1.84 8.88 2.12 ;
        RECT  8.66 1.84 8.82 3.48 ;
        RECT  7.08 2.62 7.36 3.48 ;
        RECT  4.52 1.92 4.80 2.20 ;
        RECT  4.58 1.92 4.74 3.48 ;
        RECT  2.16 1.92 2.44 2.20 ;
        RECT  2.24 1.92 2.40 3.48 ;
        RECT  0.62 1.97 0.90 2.25 ;
        RECT  0.68 1.97 0.84 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 9.60 0.28 ;
        RECT  9.14 -0.28 9.42 0.32 ;
        RECT  8.60 0.96 8.88 1.24 ;
        RECT  8.66 -0.28 8.82 1.24 ;
        RECT  7.08 0.96 7.36 1.24 ;
        RECT  7.18 -0.28 7.34 1.24 ;
        RECT  4.36 0.68 4.64 0.96 ;
        RECT  4.42 -0.28 4.58 0.96 ;
        RECT  1.64 0.68 1.92 0.96 ;
        RECT  1.70 -0.28 1.86 0.96 ;
        RECT  0.62 0.50 0.90 0.78 ;
        RECT  0.68 -0.28 0.84 0.78 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.08 0.50 0.38 0.78 ;
        RECT  0.08 1.00 1.16 1.16 ;
        RECT  0.88 0.94 1.16 1.22 ;
        RECT  0.08 0.50 0.24 2.25 ;
        RECT  0.08 1.97 0.38 2.25 ;
        RECT  1.14 0.50 1.48 0.78 ;
        RECT  1.14 1.97 1.48 2.25 ;
        RECT  1.32 0.50 1.48 2.70 ;
        RECT  1.28 2.42 1.56 2.70 ;
        RECT  2.68 0.68 3.04 0.96 ;
        RECT  1.76 1.60 3.04 1.76 ;
        RECT  1.76 1.60 1.92 2.20 ;
        RECT  1.64 1.92 1.92 2.20 ;
        RECT  2.88 0.68 3.04 2.20 ;
        RECT  2.68 1.92 3.04 2.20 ;
        RECT  3.20 0.68 3.48 0.96 ;
        RECT  3.26 0.68 3.42 2.20 ;
        RECT  3.20 1.92 3.48 2.20 ;
        RECT  3.32 1.92 3.48 2.70 ;
        RECT  3.86 2.42 4.14 2.70 ;
        RECT  3.32 2.54 4.14 2.70 ;
        RECT  3.72 0.68 4.08 0.96 ;
        RECT  3.92 0.68 4.08 2.20 ;
        RECT  3.86 1.92 4.14 2.20 ;
        RECT  4.88 0.68 5.20 0.96 ;
        RECT  4.38 1.44 5.20 1.60 ;
        RECT  4.38 1.38 4.66 1.66 ;
        RECT  5.04 0.68 5.20 2.20 ;
        RECT  5.04 1.92 5.32 2.20 ;
        RECT  5.56 0.44 7.02 0.60 ;
        RECT  6.74 0.44 7.02 0.80 ;
        RECT  5.44 0.76 5.72 1.04 ;
        RECT  5.56 0.44 5.72 2.20 ;
        RECT  5.56 1.92 5.84 2.20 ;
        RECT  6.56 0.96 6.84 1.24 ;
        RECT  6.56 1.46 7.56 1.62 ;
        RECT  7.28 1.40 7.56 1.68 ;
        RECT  6.56 0.96 6.72 2.12 ;
        RECT  6.56 1.84 6.84 2.12 ;
        RECT  5.96 0.76 6.24 1.04 ;
        RECT  7.60 0.96 7.88 1.24 ;
        RECT  7.60 1.84 7.88 2.12 ;
        RECT  6.08 0.76 6.24 2.20 ;
        RECT  6.20 1.92 6.36 2.44 ;
        RECT  7.72 0.96 7.88 2.44 ;
        RECT  6.20 2.28 8.12 2.44 ;
        RECT  7.84 2.28 8.12 2.62 ;
    END
END DFFDRBSP1V1_0

MACRO DFFDRBLDZSP8V1_0
    CLASS CORE ;
    FOREIGN DFFDRBLDZSP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 17.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 32.14  LAYER ME1  ;
        ANTENNADIFFAREA 15.73  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.76  LAYER ME1  ;
        ANTENNAMAXAREACAR 18.29  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  16.16 1.90 16.44 2.18 ;
        RECT  16.16 0.96 16.44 1.24 ;
        RECT  16.16 0.96 16.32 2.18 ;
        RECT  15.24 1.52 16.32 1.68 ;
        RECT  15.24 1.46 15.54 1.74 ;
        RECT  15.12 1.90 15.40 2.18 ;
        RECT  15.24 0.96 15.40 2.18 ;
        RECT  15.12 0.96 15.40 1.24 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 32.14  LAYER ME1  ;
        ANTENNADIFFAREA 15.73  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.76  LAYER ME1  ;
        ANTENNAMAXAREACAR 18.29  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.08 1.90 14.36 2.18 ;
        RECT  14.08 0.96 14.36 1.24 ;
        RECT  14.08 0.96 14.24 2.18 ;
        RECT  13.16 1.52 14.24 1.68 ;
        RECT  13.16 1.46 13.54 1.74 ;
        RECT  13.04 1.90 13.32 2.18 ;
        RECT  13.16 0.96 13.32 2.18 ;
        RECT  13.04 0.96 13.32 1.24 ;
        END
    END Q
    PIN LD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END LD
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 32.14  LAYER ME1  ;
        ANTENNADIFFAREA 15.54  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.76  LAYER ME1  ;
        ANTENNAMAXAREACAR 18.29  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.05 1.45 2.33 1.74 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.81 2.23 2.25 ;
        RECT  1.95 0.81 2.23 1.09 ;
        END
    END D
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.19 1.42 3.50 1.78 ;
        END
    END RB
    PIN TD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.80 1.12 6.34 1.28 ;
        RECT  5.80 1.12 6.13 1.40 ;
        END
    END TD
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.66 1.42 3.95 1.78 ;
        END
    END SEL
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.27 1.48 6.55 1.76 ;
        RECT  6.06 1.86 6.43 2.14 ;
        RECT  6.27 1.48 6.43 2.14 ;
        END
    END CK
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 17.20 0.28 ;
        RECT  16.74 -0.28 17.02 0.32 ;
        RECT  16.68 0.64 16.96 0.92 ;
        RECT  16.74 -0.28 16.90 0.92 ;
        RECT  15.64 0.64 15.92 0.92 ;
        RECT  15.70 -0.28 15.86 0.92 ;
        RECT  14.60 0.64 14.88 0.92 ;
        RECT  14.66 -0.28 14.82 0.92 ;
        RECT  13.56 0.64 13.84 0.92 ;
        RECT  13.62 -0.28 13.78 0.92 ;
        RECT  12.52 0.64 12.80 0.92 ;
        RECT  12.58 -0.28 12.74 0.92 ;
        RECT  11.52 0.96 11.80 1.24 ;
        RECT  11.62 -0.28 11.78 1.24 ;
        RECT  8.78 0.72 9.06 1.00 ;
        RECT  8.84 -0.28 9.00 1.00 ;
        RECT  6.08 0.68 6.36 0.96 ;
        RECT  6.14 -0.28 6.30 0.96 ;
        RECT  3.47 0.88 3.75 1.16 ;
        RECT  3.53 -0.28 3.69 1.16 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 17.20 3.48 ;
        RECT  16.74 2.88 17.02 3.48 ;
        RECT  16.68 2.22 16.96 2.50 ;
        RECT  16.74 2.22 16.90 3.48 ;
        RECT  15.64 2.22 15.92 2.50 ;
        RECT  15.70 2.22 15.86 3.48 ;
        RECT  14.60 2.22 14.88 2.50 ;
        RECT  14.66 2.22 14.82 3.48 ;
        RECT  13.56 2.22 13.84 2.50 ;
        RECT  13.62 2.22 13.78 3.48 ;
        RECT  12.52 1.90 12.80 2.18 ;
        RECT  12.58 1.90 12.74 3.48 ;
        RECT  11.52 1.84 11.80 2.12 ;
        RECT  11.58 1.84 11.74 3.48 ;
        RECT  8.96 1.92 9.24 2.20 ;
        RECT  9.02 1.92 9.18 3.48 ;
        RECT  7.44 2.52 7.72 3.48 ;
        RECT  3.23 2.52 3.51 3.48 ;
        RECT  2.43 1.94 2.71 2.22 ;
        RECT  2.53 1.94 2.69 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  0.91 0.81 1.19 1.09 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  1.03 0.81 1.19 2.64 ;
        RECT  1.03 2.48 2.37 2.64 ;
        RECT  2.09 2.48 2.37 2.76 ;
        RECT  1.55 0.49 2.89 0.65 ;
        RECT  2.61 0.44 2.89 0.72 ;
        RECT  1.55 0.49 1.71 1.09 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  3.99 0.88 4.27 1.16 ;
        RECT  4.11 1.26 4.43 1.54 ;
        RECT  4.11 0.88 4.27 2.22 ;
        RECT  3.99 1.94 4.27 2.22 ;
        RECT  4.52 0.68 4.80 0.96 ;
        RECT  2.43 0.88 2.71 1.16 ;
        RECT  2.43 1.00 3.03 1.16 ;
        RECT  2.87 1.00 3.03 2.22 ;
        RECT  2.87 1.94 3.23 2.22 ;
        RECT  4.64 0.68 4.80 2.14 ;
        RECT  2.87 2.06 3.83 2.22 ;
        RECT  3.67 2.06 3.83 2.54 ;
        RECT  4.52 1.86 4.68 2.54 ;
        RECT  3.67 2.38 4.68 2.54 ;
        RECT  5.48 0.68 5.84 0.96 ;
        RECT  5.48 0.68 5.64 2.14 ;
        RECT  5.48 1.86 5.84 2.14 ;
        RECT  6.60 0.68 6.97 0.96 ;
        RECT  6.81 1.16 7.20 1.44 ;
        RECT  6.81 0.68 6.97 2.14 ;
        RECT  6.68 1.86 6.97 2.14 ;
        RECT  5.04 0.68 5.32 0.96 ;
        RECT  7.16 0.72 7.52 1.00 ;
        RECT  5.10 0.68 5.26 2.14 ;
        RECT  5.04 1.86 5.32 2.14 ;
        RECT  7.36 0.72 7.52 2.20 ;
        RECT  7.13 1.92 7.52 2.20 ;
        RECT  5.16 1.86 5.32 2.46 ;
        RECT  7.13 1.92 7.29 2.46 ;
        RECT  5.16 2.30 7.29 2.46 ;
        RECT  8.24 0.72 8.54 1.00 ;
        RECT  8.24 0.72 8.40 2.20 ;
        RECT  8.20 1.92 8.48 2.20 ;
        RECT  7.68 0.72 8.04 1.00 ;
        RECT  9.04 1.48 9.32 1.76 ;
        RECT  8.64 1.60 9.32 1.76 ;
        RECT  7.68 1.92 8.04 2.20 ;
        RECT  7.88 0.72 8.04 2.52 ;
        RECT  8.64 1.60 8.80 2.52 ;
        RECT  7.88 2.36 8.80 2.52 ;
        RECT  9.30 0.72 9.64 1.00 ;
        RECT  8.56 1.16 9.64 1.32 ;
        RECT  8.56 1.16 8.84 1.44 ;
        RECT  9.48 0.72 9.64 2.20 ;
        RECT  9.48 1.92 9.76 2.20 ;
        RECT  10.38 0.76 10.80 1.04 ;
        RECT  10.52 1.92 10.80 2.20 ;
        RECT  10.64 0.76 10.80 2.76 ;
        RECT  10.64 2.48 10.92 2.76 ;
        RECT  9.98 0.44 11.46 0.60 ;
        RECT  11.18 0.44 11.46 0.80 ;
        RECT  9.86 0.76 10.14 1.04 ;
        RECT  9.98 0.44 10.14 2.20 ;
        RECT  9.98 1.92 10.28 2.20 ;
        RECT  11.00 0.96 11.28 1.24 ;
        RECT  11.00 1.46 11.94 1.62 ;
        RECT  11.66 1.40 11.94 1.68 ;
        RECT  11.00 0.96 11.16 2.12 ;
        RECT  11.00 1.84 11.28 2.12 ;
        RECT  12.04 0.96 12.32 1.24 ;
        RECT  12.04 1.84 12.32 2.12 ;
        RECT  12.13 0.96 12.29 2.70 ;
        RECT  12.13 2.42 12.42 2.70 ;
    END
END DFFDRBLDZSP8V1_0

MACRO DFFDRBLDZSP4V1_0
    CLASS CORE ;
    FOREIGN DFFDRBLDZSP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.27 1.48 6.55 1.76 ;
        RECT  6.06 1.86 6.43 2.14 ;
        RECT  6.27 1.48 6.43 2.14 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 28.63  LAYER ME1  ;
        ANTENNADIFFAREA 12.97  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.18  LAYER ME1  ;
        ANTENNAMAXAREACAR 24.25  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.20 1.46 14.54 1.74 ;
        RECT  14.08 1.90 14.36 2.18 ;
        RECT  14.20 0.96 14.36 2.18 ;
        RECT  14.08 0.96 14.36 1.24 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 28.63  LAYER ME1  ;
        ANTENNADIFFAREA 12.97  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.18  LAYER ME1  ;
        ANTENNAMAXAREACAR 24.25  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.04 1.90 13.32 2.18 ;
        RECT  13.04 0.96 13.32 1.24 ;
        RECT  13.04 0.96 13.20 2.18 ;
        RECT  12.86 1.46 13.20 1.74 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.66 1.42 3.95 1.78 ;
        END
    END SEL
    PIN TD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.80 1.12 6.34 1.28 ;
        RECT  5.80 1.12 6.13 1.40 ;
        END
    END TD
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.19 1.42 3.50 1.78 ;
        END
    END RB
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 28.63  LAYER ME1  ;
        ANTENNADIFFAREA 12.98  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.18  LAYER ME1  ;
        ANTENNAMAXAREACAR 24.25  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.05 1.45 2.33 1.74 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.81 2.23 2.25 ;
        RECT  1.95 0.81 2.23 1.09 ;
        END
    END D
    PIN LD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END LD
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 15.20 3.48 ;
        RECT  14.66 2.88 15.02 3.48 ;
        RECT  14.60 2.22 14.88 2.50 ;
        RECT  14.66 2.22 14.82 3.48 ;
        RECT  13.56 2.22 13.84 2.50 ;
        RECT  13.62 2.22 13.78 3.48 ;
        RECT  12.52 1.90 12.80 2.18 ;
        RECT  12.58 1.90 12.74 3.48 ;
        RECT  11.52 1.84 11.80 2.12 ;
        RECT  11.58 1.84 11.74 3.48 ;
        RECT  8.96 1.92 9.24 2.20 ;
        RECT  9.02 1.92 9.18 3.48 ;
        RECT  7.44 2.52 7.72 3.48 ;
        RECT  3.23 2.52 3.51 3.48 ;
        RECT  2.43 1.94 2.71 2.22 ;
        RECT  2.53 1.94 2.69 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 15.20 0.28 ;
        RECT  14.66 -0.28 15.02 0.32 ;
        RECT  14.60 0.64 14.88 0.92 ;
        RECT  14.66 -0.28 14.82 0.92 ;
        RECT  13.56 0.64 13.84 0.92 ;
        RECT  13.62 -0.28 13.78 0.92 ;
        RECT  12.52 0.64 12.80 0.92 ;
        RECT  12.58 -0.28 12.74 0.92 ;
        RECT  11.52 0.96 11.80 1.24 ;
        RECT  11.62 -0.28 11.78 1.24 ;
        RECT  8.78 0.72 9.06 1.00 ;
        RECT  8.84 -0.28 9.00 1.00 ;
        RECT  6.08 0.68 6.36 0.96 ;
        RECT  6.14 -0.28 6.30 0.96 ;
        RECT  3.47 0.88 3.75 1.16 ;
        RECT  3.53 -0.28 3.69 1.16 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  0.91 0.81 1.19 1.09 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  1.03 0.81 1.19 2.64 ;
        RECT  1.03 2.48 2.37 2.64 ;
        RECT  2.09 2.48 2.37 2.76 ;
        RECT  1.55 0.49 2.89 0.65 ;
        RECT  2.61 0.44 2.89 0.72 ;
        RECT  1.55 0.49 1.71 1.09 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  3.99 0.88 4.27 1.16 ;
        RECT  4.11 1.26 4.43 1.54 ;
        RECT  4.11 0.88 4.27 2.22 ;
        RECT  3.99 1.94 4.27 2.22 ;
        RECT  4.52 0.68 4.80 0.96 ;
        RECT  2.43 0.88 2.71 1.16 ;
        RECT  2.43 1.00 3.03 1.16 ;
        RECT  2.87 1.00 3.03 2.22 ;
        RECT  2.87 1.94 3.23 2.22 ;
        RECT  4.64 0.68 4.80 2.14 ;
        RECT  2.87 2.06 3.83 2.22 ;
        RECT  3.67 2.06 3.83 2.54 ;
        RECT  4.52 1.86 4.68 2.54 ;
        RECT  3.67 2.38 4.68 2.54 ;
        RECT  5.48 0.68 5.84 0.96 ;
        RECT  5.48 0.68 5.64 2.14 ;
        RECT  5.48 1.86 5.84 2.14 ;
        RECT  6.60 0.68 6.97 0.96 ;
        RECT  6.81 1.16 7.20 1.44 ;
        RECT  6.81 0.68 6.97 2.14 ;
        RECT  6.68 1.86 6.97 2.14 ;
        RECT  5.04 0.68 5.32 0.96 ;
        RECT  7.16 0.72 7.52 1.00 ;
        RECT  5.10 0.68 5.26 2.14 ;
        RECT  5.04 1.86 5.32 2.14 ;
        RECT  7.36 0.72 7.52 2.20 ;
        RECT  7.13 1.92 7.52 2.20 ;
        RECT  5.16 1.86 5.32 2.46 ;
        RECT  7.13 1.92 7.29 2.46 ;
        RECT  5.16 2.30 7.29 2.46 ;
        RECT  8.24 0.72 8.54 1.00 ;
        RECT  8.24 0.72 8.40 2.20 ;
        RECT  8.20 1.92 8.48 2.20 ;
        RECT  7.68 0.72 8.04 1.00 ;
        RECT  9.04 1.48 9.32 1.76 ;
        RECT  8.64 1.60 9.32 1.76 ;
        RECT  7.68 1.92 8.04 2.20 ;
        RECT  7.88 0.72 8.04 2.52 ;
        RECT  8.64 1.60 8.80 2.52 ;
        RECT  7.88 2.36 8.80 2.52 ;
        RECT  9.30 0.72 9.64 1.00 ;
        RECT  8.56 1.16 9.64 1.32 ;
        RECT  8.56 1.16 8.84 1.44 ;
        RECT  9.48 0.72 9.64 2.20 ;
        RECT  9.48 1.92 9.76 2.20 ;
        RECT  10.38 0.76 10.80 1.04 ;
        RECT  10.52 1.92 10.80 2.20 ;
        RECT  10.64 0.76 10.80 2.76 ;
        RECT  10.64 2.48 10.92 2.76 ;
        RECT  9.98 0.44 11.46 0.60 ;
        RECT  11.18 0.44 11.46 0.80 ;
        RECT  9.86 0.76 10.14 1.04 ;
        RECT  9.98 0.44 10.14 2.20 ;
        RECT  9.98 1.92 10.28 2.20 ;
        RECT  11.00 0.96 11.28 1.24 ;
        RECT  11.00 1.46 11.94 1.62 ;
        RECT  11.66 1.40 11.94 1.68 ;
        RECT  11.00 0.96 11.16 2.12 ;
        RECT  11.00 1.84 11.28 2.12 ;
        RECT  12.04 0.96 12.32 1.24 ;
        RECT  12.04 1.84 12.32 2.12 ;
        RECT  12.13 0.96 12.29 2.70 ;
        RECT  12.13 2.42 12.42 2.70 ;
    END
END DFFDRBLDZSP4V1_0

MACRO DFFDRBLDZSP2V1_0
    CLASS CORE ;
    FOREIGN DFFDRBLDZSP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN LD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END LD
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 26.67  LAYER ME1  ;
        ANTENNADIFFAREA 11.64  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.89  LAYER ME1  ;
        ANTENNAMAXAREACAR 29.87  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.05 1.45 2.33 1.74 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.81 2.23 2.25 ;
        RECT  1.95 0.81 2.23 1.09 ;
        END
    END D
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.19 1.42 3.50 1.78 ;
        END
    END RB
    PIN TD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.80 1.12 6.34 1.28 ;
        RECT  5.80 1.12 6.13 1.40 ;
        END
    END TD
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.66 1.42 3.95 1.78 ;
        END
    END SEL
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 26.67  LAYER ME1  ;
        ANTENNADIFFAREA 11.53  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.89  LAYER ME1  ;
        ANTENNAMAXAREACAR 29.87  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.52 1.90 12.80 2.18 ;
        RECT  12.52 0.96 12.80 1.24 ;
        RECT  12.52 0.96 12.74 2.18 ;
        RECT  12.46 1.46 12.74 1.74 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 26.37  LAYER ME1  ;
        ANTENNADIFFAREA 11.53  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.89  LAYER ME1  ;
        ANTENNAMAXAREACAR 29.54  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.66 1.46 13.92 1.74 ;
        RECT  13.56 1.90 13.84 2.18 ;
        RECT  13.66 0.96 13.84 2.18 ;
        RECT  13.56 0.96 13.84 1.24 ;
        END
    END QB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.27 1.48 6.55 1.76 ;
        RECT  6.06 1.86 6.43 2.14 ;
        RECT  6.27 1.48 6.43 2.14 ;
        END
    END CK
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 14.00 0.28 ;
        RECT  13.54 -0.28 13.82 0.32 ;
        RECT  13.04 0.64 13.32 0.92 ;
        RECT  13.10 -0.28 13.26 0.92 ;
        RECT  11.52 0.96 11.80 1.24 ;
        RECT  11.62 -0.28 11.78 1.24 ;
        RECT  8.78 0.72 9.06 1.00 ;
        RECT  8.84 -0.28 9.00 1.00 ;
        RECT  6.08 0.68 6.36 0.96 ;
        RECT  6.14 -0.28 6.30 0.96 ;
        RECT  3.47 0.88 3.75 1.16 ;
        RECT  3.53 -0.28 3.69 1.16 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 14.00 3.48 ;
        RECT  13.54 2.88 13.82 3.48 ;
        RECT  13.04 2.22 13.32 2.50 ;
        RECT  13.10 2.22 13.26 3.48 ;
        RECT  11.52 1.84 11.80 2.12 ;
        RECT  11.58 1.84 11.74 3.48 ;
        RECT  8.96 1.92 9.24 2.20 ;
        RECT  9.02 1.92 9.18 3.48 ;
        RECT  7.44 2.52 7.72 3.48 ;
        RECT  3.23 2.52 3.51 3.48 ;
        RECT  2.43 1.94 2.71 2.22 ;
        RECT  2.53 1.94 2.69 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  0.91 0.81 1.19 1.09 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  1.03 0.81 1.19 2.64 ;
        RECT  1.03 2.48 2.37 2.64 ;
        RECT  2.09 2.48 2.37 2.76 ;
        RECT  1.55 0.49 2.89 0.65 ;
        RECT  2.61 0.44 2.89 0.72 ;
        RECT  1.55 0.49 1.71 1.09 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  3.99 0.88 4.27 1.16 ;
        RECT  4.11 1.26 4.43 1.54 ;
        RECT  4.11 0.88 4.27 2.22 ;
        RECT  3.99 1.94 4.27 2.22 ;
        RECT  4.52 0.68 4.80 0.96 ;
        RECT  2.43 0.88 2.71 1.16 ;
        RECT  2.43 1.00 3.03 1.16 ;
        RECT  2.87 1.00 3.03 2.22 ;
        RECT  2.87 1.94 3.23 2.22 ;
        RECT  4.64 0.68 4.80 2.14 ;
        RECT  2.87 2.06 3.83 2.22 ;
        RECT  3.67 2.06 3.83 2.54 ;
        RECT  4.52 1.86 4.68 2.54 ;
        RECT  3.67 2.38 4.68 2.54 ;
        RECT  5.48 0.68 5.84 0.96 ;
        RECT  5.48 0.68 5.64 2.14 ;
        RECT  5.48 1.86 5.84 2.14 ;
        RECT  6.60 0.68 6.97 0.96 ;
        RECT  6.81 1.16 7.20 1.44 ;
        RECT  6.81 0.68 6.97 2.14 ;
        RECT  6.68 1.86 6.97 2.14 ;
        RECT  5.04 0.68 5.32 0.96 ;
        RECT  7.16 0.72 7.52 1.00 ;
        RECT  5.10 0.68 5.26 2.14 ;
        RECT  5.04 1.86 5.32 2.14 ;
        RECT  7.36 0.72 7.52 2.20 ;
        RECT  7.13 1.92 7.52 2.20 ;
        RECT  5.16 1.86 5.32 2.46 ;
        RECT  7.13 1.92 7.29 2.46 ;
        RECT  5.16 2.30 7.29 2.46 ;
        RECT  8.24 0.72 8.54 1.00 ;
        RECT  8.24 0.72 8.40 2.20 ;
        RECT  8.20 1.92 8.48 2.20 ;
        RECT  7.68 0.72 8.04 1.00 ;
        RECT  9.04 1.48 9.32 1.76 ;
        RECT  8.64 1.60 9.32 1.76 ;
        RECT  7.68 1.92 8.04 2.20 ;
        RECT  7.88 0.72 8.04 2.52 ;
        RECT  8.64 1.60 8.80 2.52 ;
        RECT  7.88 2.36 8.80 2.52 ;
        RECT  9.30 0.72 9.64 1.00 ;
        RECT  8.56 1.16 9.64 1.32 ;
        RECT  8.56 1.16 8.84 1.44 ;
        RECT  9.48 0.72 9.64 2.20 ;
        RECT  9.48 1.92 9.76 2.20 ;
        RECT  10.38 0.76 10.80 1.04 ;
        RECT  10.52 1.92 10.80 2.20 ;
        RECT  10.64 0.76 10.80 2.76 ;
        RECT  10.64 2.48 10.92 2.76 ;
        RECT  9.98 0.44 11.46 0.60 ;
        RECT  11.18 0.44 11.46 0.80 ;
        RECT  9.86 0.76 10.14 1.04 ;
        RECT  9.98 0.44 10.14 2.20 ;
        RECT  9.98 1.92 10.28 2.20 ;
        RECT  11.00 0.96 11.28 1.24 ;
        RECT  11.00 1.46 11.94 1.62 ;
        RECT  11.66 1.40 11.94 1.68 ;
        RECT  11.00 0.96 11.16 2.12 ;
        RECT  11.00 1.84 11.28 2.12 ;
        RECT  12.04 0.96 12.32 1.24 ;
        RECT  12.04 1.84 12.32 2.12 ;
        RECT  12.13 0.96 12.29 2.70 ;
        RECT  12.13 2.42 12.42 2.70 ;
    END
END DFFDRBLDZSP2V1_0

MACRO DFFDRBLDZSP1V1_0
    CLASS CORE ;
    FOREIGN DFFDRBLDZSP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 26.77  LAYER ME1  ;
        ANTENNADIFFAREA 10.95  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.74  LAYER ME1  ;
        ANTENNAMAXAREACAR 36.22  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.05 1.45 2.33 1.74 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.81 2.23 2.25 ;
        RECT  1.95 0.81 2.23 1.09 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.27 1.48 6.55 1.76 ;
        RECT  6.06 1.86 6.43 2.14 ;
        RECT  6.27 1.48 6.43 2.14 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 26.47  LAYER ME1  ;
        ANTENNADIFFAREA 10.84  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.74  LAYER ME1  ;
        ANTENNAMAXAREACAR 35.81  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.66 1.46 13.92 1.74 ;
        RECT  13.56 1.90 13.84 2.18 ;
        RECT  13.66 0.96 13.84 2.18 ;
        RECT  13.56 0.96 13.84 1.24 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 26.77  LAYER ME1  ;
        ANTENNADIFFAREA 10.84  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.74  LAYER ME1  ;
        ANTENNAMAXAREACAR 36.22  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.52 1.90 12.80 2.18 ;
        RECT  12.52 0.96 12.80 1.24 ;
        RECT  12.52 0.96 12.74 2.18 ;
        RECT  12.46 1.46 12.74 1.74 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.66 1.42 3.95 1.78 ;
        END
    END SEL
    PIN TD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.80 1.12 6.34 1.28 ;
        RECT  5.80 1.12 6.13 1.40 ;
        END
    END TD
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.19 1.42 3.50 1.78 ;
        END
    END RB
    PIN LD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END LD
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 14.00 3.48 ;
        RECT  13.54 2.88 13.82 3.48 ;
        RECT  13.04 1.90 13.32 2.18 ;
        RECT  13.10 1.90 13.26 3.48 ;
        RECT  11.52 1.84 11.80 2.12 ;
        RECT  11.58 1.84 11.74 3.48 ;
        RECT  8.96 1.92 9.24 2.20 ;
        RECT  9.02 1.92 9.18 3.48 ;
        RECT  7.44 2.52 7.72 3.48 ;
        RECT  3.23 2.52 3.51 3.48 ;
        RECT  2.43 1.94 2.71 2.22 ;
        RECT  2.53 1.94 2.69 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 14.00 0.28 ;
        RECT  13.54 -0.28 13.82 0.32 ;
        RECT  13.04 0.96 13.32 1.24 ;
        RECT  13.10 -0.28 13.26 1.24 ;
        RECT  11.52 0.96 11.80 1.24 ;
        RECT  11.62 -0.28 11.78 1.24 ;
        RECT  8.78 0.72 9.06 1.00 ;
        RECT  8.84 -0.28 9.00 1.00 ;
        RECT  6.08 0.68 6.36 0.96 ;
        RECT  6.14 -0.28 6.30 0.96 ;
        RECT  3.47 0.88 3.75 1.16 ;
        RECT  3.53 -0.28 3.69 1.16 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  0.91 0.81 1.19 1.09 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  1.03 0.81 1.19 2.64 ;
        RECT  1.03 2.48 2.37 2.64 ;
        RECT  2.09 2.48 2.37 2.76 ;
        RECT  1.55 0.49 2.89 0.65 ;
        RECT  2.61 0.44 2.89 0.72 ;
        RECT  1.55 0.49 1.71 1.09 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  3.99 0.88 4.27 1.16 ;
        RECT  4.11 1.26 4.43 1.54 ;
        RECT  4.11 0.88 4.27 2.22 ;
        RECT  3.99 1.94 4.27 2.22 ;
        RECT  4.52 0.68 4.80 0.96 ;
        RECT  2.43 0.88 2.71 1.16 ;
        RECT  2.43 1.00 3.03 1.16 ;
        RECT  2.87 1.00 3.03 2.22 ;
        RECT  2.87 1.94 3.23 2.22 ;
        RECT  4.64 0.68 4.80 2.14 ;
        RECT  2.87 2.06 3.83 2.22 ;
        RECT  3.67 2.06 3.83 2.54 ;
        RECT  4.52 1.86 4.68 2.54 ;
        RECT  3.67 2.38 4.68 2.54 ;
        RECT  5.48 0.68 5.84 0.96 ;
        RECT  5.48 0.68 5.64 2.14 ;
        RECT  5.48 1.86 5.84 2.14 ;
        RECT  6.60 0.68 6.97 0.96 ;
        RECT  6.81 1.16 7.20 1.44 ;
        RECT  6.81 0.68 6.97 2.14 ;
        RECT  6.68 1.86 6.97 2.14 ;
        RECT  5.04 0.68 5.32 0.96 ;
        RECT  7.16 0.72 7.52 1.00 ;
        RECT  5.10 0.68 5.26 2.14 ;
        RECT  5.04 1.86 5.32 2.14 ;
        RECT  7.36 0.72 7.52 2.20 ;
        RECT  7.13 1.92 7.52 2.20 ;
        RECT  5.16 1.86 5.32 2.46 ;
        RECT  7.13 1.92 7.29 2.46 ;
        RECT  5.16 2.30 7.29 2.46 ;
        RECT  8.24 0.72 8.54 1.00 ;
        RECT  8.24 0.72 8.40 2.20 ;
        RECT  8.20 1.92 8.48 2.20 ;
        RECT  7.68 0.72 8.04 1.00 ;
        RECT  9.04 1.48 9.32 1.76 ;
        RECT  8.64 1.60 9.32 1.76 ;
        RECT  7.68 1.92 8.04 2.20 ;
        RECT  7.88 0.72 8.04 2.52 ;
        RECT  8.64 1.60 8.80 2.52 ;
        RECT  7.88 2.36 8.80 2.52 ;
        RECT  9.30 0.72 9.64 1.00 ;
        RECT  8.56 1.16 9.64 1.32 ;
        RECT  8.56 1.16 8.84 1.44 ;
        RECT  9.48 0.72 9.64 2.20 ;
        RECT  9.48 1.92 9.76 2.20 ;
        RECT  10.38 0.76 10.80 1.04 ;
        RECT  10.52 1.92 10.80 2.20 ;
        RECT  10.64 0.76 10.80 2.76 ;
        RECT  10.64 2.48 10.92 2.76 ;
        RECT  9.98 0.44 11.46 0.60 ;
        RECT  11.18 0.44 11.46 0.80 ;
        RECT  9.86 0.76 10.14 1.04 ;
        RECT  9.98 0.44 10.14 2.20 ;
        RECT  9.98 1.92 10.28 2.20 ;
        RECT  11.00 0.96 11.28 1.24 ;
        RECT  11.00 1.46 11.94 1.62 ;
        RECT  11.66 1.40 11.94 1.68 ;
        RECT  11.00 0.96 11.16 2.12 ;
        RECT  11.00 1.84 11.28 2.12 ;
        RECT  12.04 0.96 12.32 1.24 ;
        RECT  12.04 1.84 12.32 2.12 ;
        RECT  12.13 0.96 12.29 2.70 ;
        RECT  12.13 2.42 12.42 2.70 ;
    END
END DFFDRBLDZSP1V1_0

MACRO DFFDRBLDSP8V1_0
    CLASS CORE ;
    FOREIGN DFFDRBLDSP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 26.98  LAYER ME1  ;
        ANTENNADIFFAREA 13.32  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.69  LAYER ME1  ;
        ANTENNAMAXAREACAR 15.97  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.49 1.90 13.77 2.18 ;
        RECT  13.49 0.96 13.77 1.24 ;
        RECT  13.49 0.96 13.65 2.18 ;
        RECT  12.46 1.52 13.65 1.68 ;
        RECT  12.46 1.46 12.74 1.74 ;
        RECT  12.45 1.90 12.73 2.18 ;
        RECT  12.46 0.96 12.73 2.18 ;
        RECT  12.45 0.96 12.73 1.24 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 26.98  LAYER ME1  ;
        ANTENNADIFFAREA 13.32  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.69  LAYER ME1  ;
        ANTENNAMAXAREACAR 15.97  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.41 1.90 11.69 2.18 ;
        RECT  11.41 0.96 11.69 1.24 ;
        RECT  11.41 0.96 11.57 2.18 ;
        RECT  10.46 1.52 11.57 1.68 ;
        RECT  10.46 1.46 10.74 1.74 ;
        RECT  10.37 1.90 10.65 2.18 ;
        RECT  10.46 0.96 10.65 2.18 ;
        RECT  10.37 0.96 10.65 1.24 ;
        END
    END Q
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.21 1.40 3.50 1.80 ;
        END
    END RB
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 26.98  LAYER ME1  ;
        ANTENNADIFFAREA 13.23  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.69  LAYER ME1  ;
        ANTENNAMAXAREACAR 15.97  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.05 1.45 2.33 1.74 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.81 2.23 2.25 ;
        RECT  1.95 0.81 2.23 1.09 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.66 1.40 3.97 1.80 ;
        END
    END CK
    PIN LD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END LD
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 14.40 0.28 ;
        RECT  14.01 0.64 14.29 0.92 ;
        RECT  14.07 -0.28 14.23 0.92 ;
        RECT  13.94 -0.28 14.23 0.32 ;
        RECT  12.97 0.64 13.25 0.92 ;
        RECT  13.03 -0.28 13.19 0.92 ;
        RECT  11.93 0.64 12.21 0.92 ;
        RECT  11.99 -0.28 12.15 0.92 ;
        RECT  10.89 0.64 11.17 0.92 ;
        RECT  10.95 -0.28 11.11 0.92 ;
        RECT  9.85 0.64 10.13 0.92 ;
        RECT  9.91 -0.28 10.07 0.92 ;
        RECT  8.85 0.96 9.13 1.24 ;
        RECT  8.95 -0.28 9.11 1.24 ;
        RECT  6.11 0.72 6.39 1.00 ;
        RECT  6.17 -0.28 6.33 1.00 ;
        RECT  3.47 0.88 3.75 1.16 ;
        RECT  3.53 -0.28 3.69 1.16 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 14.40 3.48 ;
        RECT  14.01 2.22 14.29 2.50 ;
        RECT  13.94 2.88 14.23 3.48 ;
        RECT  14.07 2.22 14.23 3.48 ;
        RECT  12.97 2.22 13.25 2.50 ;
        RECT  13.03 2.22 13.19 3.48 ;
        RECT  11.93 2.22 12.21 2.50 ;
        RECT  11.99 2.22 12.15 3.48 ;
        RECT  10.89 2.22 11.17 2.50 ;
        RECT  10.95 2.22 11.11 3.48 ;
        RECT  9.85 1.90 10.13 2.18 ;
        RECT  9.91 1.90 10.07 3.48 ;
        RECT  8.85 1.84 9.13 2.12 ;
        RECT  8.91 1.84 9.07 3.48 ;
        RECT  6.29 1.92 6.57 2.20 ;
        RECT  6.35 1.92 6.51 3.48 ;
        RECT  3.25 2.52 3.53 3.48 ;
        RECT  2.43 1.96 2.71 2.24 ;
        RECT  2.53 1.96 2.69 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  0.91 0.81 1.19 1.09 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  1.03 0.81 1.19 2.64 ;
        RECT  1.03 2.48 2.37 2.64 ;
        RECT  2.09 2.48 2.37 2.76 ;
        RECT  1.55 0.49 2.90 0.65 ;
        RECT  2.62 0.44 2.90 0.72 ;
        RECT  1.55 0.49 1.71 1.09 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  3.99 0.88 4.33 1.16 ;
        RECT  4.17 1.26 4.45 1.54 ;
        RECT  4.17 0.88 4.33 2.24 ;
        RECT  4.01 1.96 4.33 2.24 ;
        RECT  2.43 0.88 2.71 1.16 ;
        RECT  4.49 0.72 4.77 1.00 ;
        RECT  2.43 1.00 3.03 1.16 ;
        RECT  2.87 1.00 3.03 2.24 ;
        RECT  2.87 1.96 3.23 2.24 ;
        RECT  4.61 0.72 4.77 2.20 ;
        RECT  2.87 2.08 3.85 2.24 ;
        RECT  3.69 2.08 3.85 2.56 ;
        RECT  4.49 1.92 4.65 2.56 ;
        RECT  3.69 2.40 4.65 2.56 ;
        RECT  5.57 0.72 5.87 1.00 ;
        RECT  5.57 0.72 5.73 2.20 ;
        RECT  5.53 1.92 5.81 2.20 ;
        RECT  5.01 0.72 5.29 1.00 ;
        RECT  6.37 1.48 6.65 1.76 ;
        RECT  5.97 1.60 6.65 1.76 ;
        RECT  5.07 0.72 5.23 2.20 ;
        RECT  5.01 1.92 5.29 2.20 ;
        RECT  5.13 1.92 5.29 2.52 ;
        RECT  5.97 1.60 6.13 2.52 ;
        RECT  5.13 2.36 6.13 2.52 ;
        RECT  6.63 0.72 6.97 1.00 ;
        RECT  5.89 1.16 6.97 1.32 ;
        RECT  5.89 1.16 6.17 1.44 ;
        RECT  6.81 0.72 6.97 2.20 ;
        RECT  6.81 1.92 7.09 2.20 ;
        RECT  7.71 0.76 8.01 1.04 ;
        RECT  7.85 0.76 8.01 2.20 ;
        RECT  7.97 1.92 8.13 2.76 ;
        RECT  7.97 2.48 8.25 2.76 ;
        RECT  7.31 0.44 8.79 0.60 ;
        RECT  8.51 0.44 8.79 0.80 ;
        RECT  7.19 0.76 7.47 1.04 ;
        RECT  7.31 0.44 7.47 2.20 ;
        RECT  7.31 1.92 7.61 2.20 ;
        RECT  8.33 0.96 8.61 1.24 ;
        RECT  8.33 1.46 9.27 1.62 ;
        RECT  8.99 1.40 9.27 1.68 ;
        RECT  8.33 0.96 8.49 2.12 ;
        RECT  8.33 1.84 8.61 2.12 ;
        RECT  9.37 0.96 9.65 1.24 ;
        RECT  9.37 1.84 9.65 2.12 ;
        RECT  9.46 0.96 9.62 2.70 ;
        RECT  9.46 2.42 9.75 2.70 ;
    END
END DFFDRBLDSP8V1_0

MACRO DFFDRBLDSP4V1_0
    CLASS CORE ;
    FOREIGN DFFDRBLDSP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN LD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END LD
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 23.39  LAYER ME1  ;
        ANTENNADIFFAREA 10.56  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.11  LAYER ME1  ;
        ANTENNAMAXAREACAR 21.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.46 1.46 10.74 1.74 ;
        RECT  10.37 1.90 10.65 2.18 ;
        RECT  10.46 0.96 10.65 2.18 ;
        RECT  10.37 0.96 10.65 1.24 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 23.08  LAYER ME1  ;
        ANTENNADIFFAREA 10.56  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.11  LAYER ME1  ;
        ANTENNAMAXAREACAR 20.73  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.41 1.90 11.69 2.18 ;
        RECT  11.41 0.96 11.69 1.24 ;
        RECT  11.41 0.96 11.57 2.18 ;
        RECT  11.26 1.46 11.57 1.74 ;
        END
    END QB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.66 1.40 3.97 1.80 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 23.39  LAYER ME1  ;
        ANTENNADIFFAREA 10.67  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.11  LAYER ME1  ;
        ANTENNAMAXAREACAR 21.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.05 1.45 2.33 1.74 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.81 2.23 2.25 ;
        RECT  1.95 0.81 2.23 1.09 ;
        END
    END D
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.21 1.40 3.50 1.80 ;
        END
    END RB
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 12.40 0.28 ;
        RECT  11.94 -0.28 12.22 0.32 ;
        RECT  11.93 0.64 12.21 0.92 ;
        RECT  11.99 -0.28 12.15 0.92 ;
        RECT  10.89 0.64 11.17 0.92 ;
        RECT  10.95 -0.28 11.11 0.92 ;
        RECT  9.85 0.64 10.13 0.92 ;
        RECT  9.91 -0.28 10.07 0.92 ;
        RECT  8.85 0.96 9.13 1.24 ;
        RECT  8.95 -0.28 9.11 1.24 ;
        RECT  6.11 0.72 6.39 1.00 ;
        RECT  6.17 -0.28 6.33 1.00 ;
        RECT  3.47 0.88 3.75 1.16 ;
        RECT  3.53 -0.28 3.69 1.16 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 12.40 3.48 ;
        RECT  11.94 2.88 12.22 3.48 ;
        RECT  11.93 2.22 12.21 2.50 ;
        RECT  11.99 2.22 12.15 3.48 ;
        RECT  10.89 2.22 11.17 2.50 ;
        RECT  10.95 2.22 11.11 3.48 ;
        RECT  9.85 1.90 10.13 2.18 ;
        RECT  9.91 1.90 10.07 3.48 ;
        RECT  8.85 1.84 9.13 2.12 ;
        RECT  8.91 1.84 9.07 3.48 ;
        RECT  6.29 1.92 6.57 2.20 ;
        RECT  6.35 1.92 6.51 3.48 ;
        RECT  3.25 2.52 3.53 3.48 ;
        RECT  2.43 1.96 2.71 2.24 ;
        RECT  2.53 1.96 2.69 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  0.91 0.81 1.19 1.09 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  1.03 0.81 1.19 2.64 ;
        RECT  1.03 2.48 2.37 2.64 ;
        RECT  2.09 2.48 2.37 2.76 ;
        RECT  1.55 0.49 2.90 0.65 ;
        RECT  2.62 0.44 2.90 0.72 ;
        RECT  1.55 0.49 1.71 1.09 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  3.99 0.88 4.33 1.16 ;
        RECT  4.17 1.26 4.45 1.54 ;
        RECT  4.17 0.88 4.33 2.24 ;
        RECT  4.01 1.96 4.33 2.24 ;
        RECT  2.43 0.88 2.71 1.16 ;
        RECT  4.49 0.72 4.77 1.00 ;
        RECT  2.43 1.00 3.03 1.16 ;
        RECT  2.87 1.00 3.03 2.24 ;
        RECT  2.87 1.96 3.23 2.24 ;
        RECT  4.61 0.72 4.77 2.20 ;
        RECT  2.87 2.08 3.85 2.24 ;
        RECT  3.69 2.08 3.85 2.56 ;
        RECT  4.49 1.92 4.65 2.56 ;
        RECT  3.69 2.40 4.65 2.56 ;
        RECT  5.57 0.72 5.87 1.00 ;
        RECT  5.57 0.72 5.73 2.20 ;
        RECT  5.53 1.92 5.81 2.20 ;
        RECT  5.01 0.72 5.29 1.00 ;
        RECT  6.37 1.48 6.65 1.76 ;
        RECT  5.97 1.60 6.65 1.76 ;
        RECT  5.07 0.72 5.23 2.20 ;
        RECT  5.01 1.92 5.29 2.20 ;
        RECT  5.13 1.92 5.29 2.52 ;
        RECT  5.97 1.60 6.13 2.52 ;
        RECT  5.13 2.36 6.13 2.52 ;
        RECT  6.63 0.72 6.97 1.00 ;
        RECT  5.89 1.16 6.97 1.32 ;
        RECT  5.89 1.16 6.17 1.44 ;
        RECT  6.81 0.72 6.97 2.20 ;
        RECT  6.81 1.92 7.09 2.20 ;
        RECT  7.71 0.76 8.01 1.04 ;
        RECT  7.85 0.76 8.01 2.20 ;
        RECT  7.97 1.92 8.13 2.76 ;
        RECT  7.97 2.48 8.25 2.76 ;
        RECT  7.31 0.44 8.79 0.60 ;
        RECT  8.51 0.44 8.79 0.80 ;
        RECT  7.19 0.76 7.47 1.04 ;
        RECT  7.31 0.44 7.47 2.20 ;
        RECT  7.31 1.92 7.61 2.20 ;
        RECT  8.33 0.96 8.61 1.24 ;
        RECT  8.33 1.46 9.27 1.62 ;
        RECT  8.99 1.40 9.27 1.68 ;
        RECT  8.33 0.96 8.49 2.12 ;
        RECT  8.33 1.84 8.61 2.12 ;
        RECT  9.37 0.96 9.65 1.24 ;
        RECT  9.37 1.84 9.65 2.12 ;
        RECT  9.46 0.96 9.62 2.70 ;
        RECT  9.46 2.42 9.75 2.70 ;
    END
END DFFDRBLDSP4V1_0

MACRO DFFDRBLDSP2V1_0
    CLASS CORE ;
    FOREIGN DFFDRBLDSP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.21 1.40 3.50 1.80 ;
        END
    END RB
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 21.93  LAYER ME1  ;
        ANTENNADIFFAREA 9.45  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.83  LAYER ME1  ;
        ANTENNAMAXAREACAR 26.56  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.05 1.45 2.33 1.74 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.81 2.23 2.25 ;
        RECT  1.95 0.81 2.23 1.09 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.66 1.40 3.97 1.80 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 21.93  LAYER ME1  ;
        ANTENNADIFFAREA 9.34  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.83  LAYER ME1  ;
        ANTENNAMAXAREACAR 26.56  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.89 1.90 11.17 2.18 ;
        RECT  10.89 0.96 11.17 1.24 ;
        RECT  10.89 0.96 11.14 2.18 ;
        RECT  10.86 1.46 11.14 1.74 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 21.93  LAYER ME1  ;
        ANTENNADIFFAREA 9.34  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.83  LAYER ME1  ;
        ANTENNAMAXAREACAR 26.56  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.97 1.46 10.34 1.74 ;
        RECT  9.85 1.90 10.13 2.18 ;
        RECT  9.97 0.96 10.13 2.18 ;
        RECT  9.85 0.96 10.13 1.24 ;
        END
    END Q
    PIN LD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END LD
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 11.60 3.48 ;
        RECT  11.14 2.88 11.42 3.48 ;
        RECT  10.37 2.22 10.65 2.50 ;
        RECT  10.43 2.22 10.59 3.48 ;
        RECT  8.85 1.84 9.13 2.12 ;
        RECT  8.91 1.84 9.07 3.48 ;
        RECT  6.29 1.92 6.57 2.20 ;
        RECT  6.35 1.92 6.51 3.48 ;
        RECT  3.25 2.52 3.53 3.48 ;
        RECT  2.43 1.96 2.71 2.24 ;
        RECT  2.53 1.96 2.69 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 11.60 0.28 ;
        RECT  11.14 -0.28 11.42 0.32 ;
        RECT  10.37 0.64 10.65 0.92 ;
        RECT  10.43 -0.28 10.59 0.92 ;
        RECT  8.85 0.96 9.13 1.24 ;
        RECT  8.95 -0.28 9.11 1.24 ;
        RECT  6.11 0.72 6.39 1.00 ;
        RECT  6.17 -0.28 6.33 1.00 ;
        RECT  3.47 0.88 3.75 1.16 ;
        RECT  3.53 -0.28 3.69 1.16 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  0.91 0.81 1.19 1.09 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  1.03 0.81 1.19 2.64 ;
        RECT  1.03 2.48 2.37 2.64 ;
        RECT  2.09 2.48 2.37 2.76 ;
        RECT  1.55 0.49 2.90 0.65 ;
        RECT  2.62 0.44 2.90 0.72 ;
        RECT  1.55 0.49 1.71 1.09 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  3.99 0.88 4.33 1.16 ;
        RECT  4.17 1.26 4.45 1.54 ;
        RECT  4.17 0.88 4.33 2.24 ;
        RECT  4.01 1.96 4.33 2.24 ;
        RECT  2.43 0.88 2.71 1.16 ;
        RECT  4.49 0.72 4.77 1.00 ;
        RECT  2.43 1.00 3.03 1.16 ;
        RECT  2.87 1.00 3.03 2.24 ;
        RECT  2.87 1.96 3.23 2.24 ;
        RECT  4.61 0.72 4.77 2.20 ;
        RECT  2.87 2.08 3.85 2.24 ;
        RECT  3.69 2.08 3.85 2.56 ;
        RECT  4.49 1.92 4.65 2.56 ;
        RECT  3.69 2.40 4.65 2.56 ;
        RECT  5.57 0.72 5.87 1.00 ;
        RECT  5.57 0.72 5.73 2.20 ;
        RECT  5.53 1.92 5.81 2.20 ;
        RECT  5.01 0.72 5.29 1.00 ;
        RECT  6.37 1.48 6.65 1.76 ;
        RECT  5.97 1.60 6.65 1.76 ;
        RECT  5.07 0.72 5.23 2.20 ;
        RECT  5.01 1.92 5.29 2.20 ;
        RECT  5.13 1.92 5.29 2.52 ;
        RECT  5.97 1.60 6.13 2.52 ;
        RECT  5.13 2.36 6.13 2.52 ;
        RECT  6.63 0.72 6.97 1.00 ;
        RECT  5.89 1.16 6.97 1.32 ;
        RECT  5.89 1.16 6.17 1.44 ;
        RECT  6.81 0.72 6.97 2.20 ;
        RECT  6.81 1.92 7.09 2.20 ;
        RECT  7.71 0.76 8.01 1.04 ;
        RECT  7.85 0.76 8.01 2.20 ;
        RECT  7.97 1.92 8.13 2.76 ;
        RECT  7.97 2.48 8.25 2.76 ;
        RECT  7.31 0.44 8.79 0.60 ;
        RECT  8.51 0.44 8.79 0.80 ;
        RECT  7.19 0.76 7.47 1.04 ;
        RECT  7.31 0.44 7.47 2.20 ;
        RECT  7.31 1.92 7.61 2.20 ;
        RECT  8.33 0.96 8.61 1.24 ;
        RECT  8.33 1.46 9.27 1.62 ;
        RECT  8.99 1.40 9.27 1.68 ;
        RECT  8.33 0.96 8.49 2.12 ;
        RECT  8.33 1.84 8.61 2.12 ;
        RECT  9.37 0.96 9.65 1.24 ;
        RECT  9.37 1.84 9.65 2.12 ;
        RECT  9.46 0.96 9.62 2.70 ;
        RECT  9.46 2.42 9.75 2.70 ;
    END
END DFFDRBLDSP2V1_0

MACRO DFFDRBLDSP1V1_0
    CLASS CORE ;
    FOREIGN DFFDRBLDSP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 22.03  LAYER ME1  ;
        ANTENNADIFFAREA 8.65  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER ME1  ;
        ANTENNAMAXAREACAR 32.79  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.97 1.46 10.34 1.74 ;
        RECT  9.85 1.90 10.13 2.18 ;
        RECT  9.97 0.96 10.13 2.18 ;
        RECT  9.85 0.96 10.13 1.24 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 22.03  LAYER ME1  ;
        ANTENNADIFFAREA 8.65  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER ME1  ;
        ANTENNAMAXAREACAR 32.79  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.89 1.90 11.17 2.18 ;
        RECT  10.89 0.96 11.17 1.24 ;
        RECT  10.89 0.96 11.14 2.18 ;
        RECT  10.86 1.46 11.14 1.74 ;
        END
    END QB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.66 1.40 3.97 1.80 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 22.03  LAYER ME1  ;
        ANTENNADIFFAREA 8.76  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER ME1  ;
        ANTENNAMAXAREACAR 32.79  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.05 1.45 2.33 1.74 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.81 2.23 2.25 ;
        RECT  1.95 0.81 2.23 1.09 ;
        END
    END D
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.21 1.40 3.50 1.80 ;
        END
    END RB
    PIN LD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END LD
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 11.60 0.28 ;
        RECT  11.14 -0.28 11.42 0.32 ;
        RECT  10.37 0.96 10.65 1.24 ;
        RECT  10.43 -0.28 10.59 1.24 ;
        RECT  8.85 0.96 9.13 1.24 ;
        RECT  8.95 -0.28 9.11 1.24 ;
        RECT  6.11 0.72 6.39 1.00 ;
        RECT  6.17 -0.28 6.33 1.00 ;
        RECT  3.47 0.88 3.75 1.16 ;
        RECT  3.53 -0.28 3.69 1.16 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 11.60 3.48 ;
        RECT  11.14 2.88 11.42 3.48 ;
        RECT  10.37 1.90 10.65 2.18 ;
        RECT  10.43 1.90 10.59 3.48 ;
        RECT  8.85 1.84 9.13 2.12 ;
        RECT  8.91 1.84 9.07 3.48 ;
        RECT  6.29 1.92 6.57 2.20 ;
        RECT  6.35 1.92 6.51 3.48 ;
        RECT  3.25 2.52 3.53 3.48 ;
        RECT  2.43 1.96 2.71 2.24 ;
        RECT  2.53 1.96 2.69 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  0.91 0.81 1.19 1.09 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  1.03 0.81 1.19 2.64 ;
        RECT  1.03 2.48 2.37 2.64 ;
        RECT  2.09 2.48 2.37 2.76 ;
        RECT  1.55 0.49 2.90 0.65 ;
        RECT  2.62 0.44 2.90 0.72 ;
        RECT  1.55 0.49 1.71 1.09 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  3.99 0.88 4.33 1.16 ;
        RECT  4.17 1.26 4.45 1.54 ;
        RECT  4.17 0.88 4.33 2.24 ;
        RECT  4.01 1.96 4.33 2.24 ;
        RECT  2.43 0.88 2.71 1.16 ;
        RECT  4.49 0.72 4.77 1.00 ;
        RECT  2.43 1.00 3.03 1.16 ;
        RECT  2.87 1.00 3.03 2.24 ;
        RECT  2.87 1.96 3.23 2.24 ;
        RECT  4.61 0.72 4.77 2.20 ;
        RECT  2.87 2.08 3.85 2.24 ;
        RECT  3.69 2.08 3.85 2.56 ;
        RECT  4.49 1.92 4.65 2.56 ;
        RECT  3.69 2.40 4.65 2.56 ;
        RECT  5.57 0.72 5.87 1.00 ;
        RECT  5.57 0.72 5.73 2.20 ;
        RECT  5.53 1.92 5.81 2.20 ;
        RECT  5.01 0.72 5.29 1.00 ;
        RECT  6.37 1.48 6.65 1.76 ;
        RECT  5.97 1.60 6.65 1.76 ;
        RECT  5.07 0.72 5.23 2.20 ;
        RECT  5.01 1.92 5.29 2.20 ;
        RECT  5.13 1.92 5.29 2.52 ;
        RECT  5.97 1.60 6.13 2.52 ;
        RECT  5.13 2.36 6.13 2.52 ;
        RECT  6.63 0.72 6.97 1.00 ;
        RECT  5.89 1.16 6.97 1.32 ;
        RECT  5.89 1.16 6.17 1.44 ;
        RECT  6.81 0.72 6.97 2.20 ;
        RECT  6.81 1.92 7.09 2.20 ;
        RECT  7.71 0.76 8.01 1.04 ;
        RECT  7.85 0.76 8.01 2.20 ;
        RECT  7.97 1.92 8.13 2.76 ;
        RECT  7.97 2.48 8.25 2.76 ;
        RECT  7.31 0.44 8.79 0.60 ;
        RECT  8.51 0.44 8.79 0.80 ;
        RECT  7.19 0.76 7.47 1.04 ;
        RECT  7.31 0.44 7.47 2.20 ;
        RECT  7.31 1.92 7.61 2.20 ;
        RECT  8.33 0.96 8.61 1.24 ;
        RECT  8.33 1.46 9.27 1.62 ;
        RECT  8.99 1.40 9.27 1.68 ;
        RECT  8.33 0.96 8.49 2.12 ;
        RECT  8.33 1.84 8.61 2.12 ;
        RECT  9.37 0.96 9.65 1.24 ;
        RECT  9.37 1.84 9.65 2.12 ;
        RECT  9.46 0.96 9.62 2.70 ;
        RECT  9.46 2.42 9.75 2.70 ;
    END
END DFFDRBLDSP1V1_0

MACRO DFFDEZSP8V1_0
    CLASS CORE ;
    FOREIGN DFFDEZSP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 30.58  LAYER ME1  ;
        ANTENNADIFFAREA 14.95  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.76  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.41  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  15.32 1.90 15.60 2.18 ;
        RECT  15.32 0.96 15.60 1.24 ;
        RECT  15.32 0.96 15.48 2.18 ;
        RECT  14.40 1.52 15.48 1.68 ;
        RECT  14.40 1.46 14.74 1.74 ;
        RECT  14.28 1.90 14.56 2.18 ;
        RECT  14.40 0.96 14.56 2.18 ;
        RECT  14.28 0.96 14.56 1.24 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 30.58  LAYER ME1  ;
        ANTENNADIFFAREA 14.86  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.76  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.41  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.21 1.88 1.51 2.16 ;
        RECT  1.21 0.66 1.51 0.96 ;
        RECT  1.21 0.66 1.37 2.16 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.99 1.46 2.34 1.76 ;
        END
    END E
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.45 1.06 2.78 1.34 ;
        RECT  2.26 1.06 2.78 1.30 ;
        END
    END SEL
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 30.58  LAYER ME1  ;
        ANTENNADIFFAREA 14.95  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.76  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.41  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.24 1.90 13.52 2.18 ;
        RECT  13.24 0.96 13.52 1.24 ;
        RECT  13.24 0.96 13.40 2.18 ;
        RECT  12.32 1.52 13.40 1.68 ;
        RECT  12.32 1.46 12.74 1.74 ;
        RECT  12.20 1.90 12.48 2.18 ;
        RECT  12.32 0.96 12.48 2.18 ;
        RECT  12.20 0.96 12.48 1.24 ;
        END
    END Q
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.26 1.46 5.72 1.74 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 30.58  LAYER ME1  ;
        ANTENNADIFFAREA 14.86  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.76  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.41  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.30 1.98 4.58 2.26 ;
        RECT  4.30 0.76 4.58 1.04 ;
        RECT  4.30 0.76 4.46 2.26 ;
        RECT  4.06 1.46 4.46 1.74 ;
        END
    END TD
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 16.40 0.28 ;
        RECT  15.90 -0.28 16.22 0.32 ;
        RECT  15.84 0.64 16.12 0.92 ;
        RECT  15.90 -0.28 16.06 0.92 ;
        RECT  14.80 0.64 15.08 0.92 ;
        RECT  14.86 -0.28 15.02 0.92 ;
        RECT  13.76 0.64 14.04 0.92 ;
        RECT  13.82 -0.28 13.98 0.92 ;
        RECT  12.72 0.64 13.00 0.92 ;
        RECT  12.78 -0.28 12.94 0.92 ;
        RECT  11.68 0.64 11.96 0.92 ;
        RECT  11.74 -0.28 11.90 0.92 ;
        RECT  10.68 0.96 10.96 1.24 ;
        RECT  10.78 -0.28 10.94 1.24 ;
        RECT  7.94 0.72 8.22 1.00 ;
        RECT  8.00 -0.28 8.16 1.00 ;
        RECT  5.30 0.88 5.58 1.16 ;
        RECT  5.40 -0.28 5.56 1.16 ;
        RECT  2.26 0.62 2.54 0.90 ;
        RECT  2.32 -0.28 2.48 0.90 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 16.40 3.48 ;
        RECT  15.90 2.88 16.22 3.48 ;
        RECT  15.84 2.22 16.12 2.50 ;
        RECT  15.90 2.22 16.06 3.48 ;
        RECT  14.80 2.22 15.08 2.50 ;
        RECT  14.86 2.22 15.02 3.48 ;
        RECT  13.76 2.22 14.04 2.50 ;
        RECT  13.82 2.22 13.98 3.48 ;
        RECT  12.72 2.22 13.00 2.50 ;
        RECT  12.78 2.22 12.94 3.48 ;
        RECT  11.68 2.22 11.96 2.50 ;
        RECT  11.74 2.22 11.90 3.48 ;
        RECT  10.68 1.84 10.96 2.12 ;
        RECT  10.74 1.84 10.90 3.48 ;
        RECT  8.12 1.92 8.40 2.20 ;
        RECT  8.18 1.92 8.34 3.48 ;
        RECT  5.09 2.52 5.37 3.48 ;
        RECT  3.78 2.52 4.06 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.19 0.68 0.47 0.96 ;
        RECT  0.19 1.88 0.47 2.16 ;
        RECT  0.19 0.68 0.35 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  1.67 0.62 2.02 0.90 ;
        RECT  1.53 1.12 1.83 1.40 ;
        RECT  1.67 0.62 1.83 2.20 ;
        RECT  1.67 1.92 2.02 2.20 ;
        RECT  2.78 0.62 3.10 0.90 ;
        RECT  2.94 1.22 3.22 1.50 ;
        RECT  2.94 0.62 3.10 2.20 ;
        RECT  2.78 1.92 3.10 2.20 ;
        RECT  0.71 0.68 0.99 0.96 ;
        RECT  3.26 0.76 3.54 1.04 ;
        RECT  0.77 0.68 0.93 2.16 ;
        RECT  0.71 1.88 0.99 2.16 ;
        RECT  3.38 0.76 3.54 2.26 ;
        RECT  0.83 1.88 0.99 2.52 ;
        RECT  3.26 1.98 3.42 2.52 ;
        RECT  0.83 2.36 3.42 2.52 ;
        RECT  3.90 0.44 5.24 0.60 ;
        RECT  4.96 0.44 5.24 0.72 ;
        RECT  3.90 0.44 4.06 1.04 ;
        RECT  3.74 0.76 3.90 2.26 ;
        RECT  3.74 1.98 4.06 2.26 ;
        RECT  5.82 0.88 6.12 1.16 ;
        RECT  5.96 1.26 6.24 1.54 ;
        RECT  5.96 0.88 6.12 2.14 ;
        RECT  5.84 1.86 6.12 2.14 ;
        RECT  6.32 0.72 6.60 1.00 ;
        RECT  4.78 0.88 5.06 1.16 ;
        RECT  4.78 0.88 4.94 2.14 ;
        RECT  6.40 0.72 6.56 2.20 ;
        RECT  4.78 1.86 5.06 2.14 ;
        RECT  4.78 1.98 5.68 2.14 ;
        RECT  6.32 1.92 6.60 2.20 ;
        RECT  5.52 1.98 5.68 2.46 ;
        RECT  6.32 1.92 6.48 2.46 ;
        RECT  5.52 2.30 6.48 2.46 ;
        RECT  7.40 0.72 7.70 1.00 ;
        RECT  7.40 0.72 7.56 2.20 ;
        RECT  7.36 1.92 7.64 2.20 ;
        RECT  6.84 0.72 7.12 1.00 ;
        RECT  8.20 1.48 8.48 1.76 ;
        RECT  7.80 1.60 8.48 1.76 ;
        RECT  6.90 0.72 7.06 2.20 ;
        RECT  6.84 1.92 7.12 2.20 ;
        RECT  6.96 1.92 7.12 2.52 ;
        RECT  7.80 1.60 7.96 2.52 ;
        RECT  6.96 2.36 7.96 2.52 ;
        RECT  8.46 0.72 8.80 1.00 ;
        RECT  7.72 1.16 8.80 1.32 ;
        RECT  7.72 1.16 8.00 1.44 ;
        RECT  8.64 0.72 8.80 2.20 ;
        RECT  8.64 1.92 8.92 2.20 ;
        RECT  9.54 0.76 9.96 1.04 ;
        RECT  9.68 1.92 9.96 2.20 ;
        RECT  9.80 0.76 9.96 2.76 ;
        RECT  9.80 2.48 10.08 2.76 ;
        RECT  9.14 0.44 10.62 0.60 ;
        RECT  10.34 0.44 10.62 0.80 ;
        RECT  9.02 0.76 9.30 1.04 ;
        RECT  9.14 0.44 9.30 2.20 ;
        RECT  9.14 1.92 9.44 2.20 ;
        RECT  10.16 0.96 10.44 1.24 ;
        RECT  10.16 1.46 11.10 1.62 ;
        RECT  10.82 1.40 11.10 1.68 ;
        RECT  10.16 0.96 10.32 2.12 ;
        RECT  10.16 1.84 10.44 2.12 ;
        RECT  11.20 0.96 11.48 1.24 ;
        RECT  11.20 1.84 11.48 2.12 ;
        RECT  11.29 0.96 11.45 2.76 ;
        RECT  11.23 2.48 11.51 2.76 ;
    END
END DFFDEZSP8V1_0

MACRO DFFDEZSP4V1_0
    CLASS CORE ;
    FOREIGN DFFDEZSP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 27.07  LAYER ME1  ;
        ANTENNADIFFAREA 12.30  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.18  LAYER ME1  ;
        ANTENNAMAXAREACAR 22.93  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.30 1.98 4.58 2.26 ;
        RECT  4.30 0.76 4.58 1.04 ;
        RECT  4.30 0.76 4.46 2.26 ;
        RECT  4.06 1.46 4.46 1.74 ;
        END
    END TD
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.26 1.46 5.72 1.74 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 26.77  LAYER ME1  ;
        ANTENNADIFFAREA 12.19  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.18  LAYER ME1  ;
        ANTENNAMAXAREACAR 22.67  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.20 1.90 12.48 2.18 ;
        RECT  12.20 0.96 12.48 1.24 ;
        RECT  12.20 0.96 12.36 2.18 ;
        RECT  12.06 1.46 12.36 1.74 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.45 1.06 2.78 1.34 ;
        RECT  2.26 1.06 2.78 1.30 ;
        END
    END SEL
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.99 1.46 2.34 1.76 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 27.07  LAYER ME1  ;
        ANTENNADIFFAREA 12.30  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.18  LAYER ME1  ;
        ANTENNAMAXAREACAR 22.93  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.21 1.88 1.51 2.16 ;
        RECT  1.21 0.66 1.51 0.96 ;
        RECT  1.21 0.66 1.37 2.16 ;
        END
    END D
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 27.07  LAYER ME1  ;
        ANTENNADIFFAREA 12.19  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.18  LAYER ME1  ;
        ANTENNAMAXAREACAR 22.93  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.26 1.46 13.54 1.74 ;
        RECT  13.24 1.90 13.52 2.18 ;
        RECT  13.26 0.96 13.52 2.18 ;
        RECT  13.24 0.96 13.52 1.24 ;
        END
    END QB
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 14.40 3.48 ;
        RECT  13.82 2.88 14.22 3.48 ;
        RECT  13.76 2.22 14.04 2.50 ;
        RECT  13.82 2.22 13.98 3.48 ;
        RECT  12.72 2.22 13.00 2.50 ;
        RECT  12.78 2.22 12.94 3.48 ;
        RECT  11.68 2.22 11.96 2.50 ;
        RECT  11.74 2.22 11.90 3.48 ;
        RECT  10.68 1.84 10.96 2.12 ;
        RECT  10.74 1.84 10.90 3.48 ;
        RECT  8.12 1.92 8.40 2.20 ;
        RECT  8.18 1.92 8.34 3.48 ;
        RECT  5.09 2.52 5.37 3.48 ;
        RECT  3.78 2.52 4.06 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 14.40 0.28 ;
        RECT  13.82 -0.28 14.22 0.32 ;
        RECT  13.76 0.64 14.04 0.92 ;
        RECT  13.82 -0.28 13.98 0.92 ;
        RECT  12.72 0.64 13.00 0.92 ;
        RECT  12.78 -0.28 12.94 0.92 ;
        RECT  11.68 0.64 11.96 0.92 ;
        RECT  11.74 -0.28 11.90 0.92 ;
        RECT  10.68 0.96 10.96 1.24 ;
        RECT  10.78 -0.28 10.94 1.24 ;
        RECT  7.94 0.72 8.22 1.00 ;
        RECT  8.00 -0.28 8.16 1.00 ;
        RECT  5.30 0.88 5.58 1.16 ;
        RECT  5.40 -0.28 5.56 1.16 ;
        RECT  2.26 0.62 2.54 0.90 ;
        RECT  2.32 -0.28 2.48 0.90 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.19 0.68 0.47 0.96 ;
        RECT  0.19 1.88 0.47 2.16 ;
        RECT  0.19 0.68 0.35 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  1.67 0.62 2.02 0.90 ;
        RECT  1.53 1.12 1.83 1.40 ;
        RECT  1.67 0.62 1.83 2.20 ;
        RECT  1.67 1.92 2.02 2.20 ;
        RECT  2.78 0.62 3.10 0.90 ;
        RECT  2.94 1.22 3.22 1.50 ;
        RECT  2.94 0.62 3.10 2.20 ;
        RECT  2.78 1.92 3.10 2.20 ;
        RECT  0.71 0.68 0.99 0.96 ;
        RECT  3.26 0.76 3.54 1.04 ;
        RECT  0.77 0.68 0.93 2.16 ;
        RECT  0.71 1.88 0.99 2.16 ;
        RECT  3.38 0.76 3.54 2.26 ;
        RECT  0.83 1.88 0.99 2.52 ;
        RECT  3.26 1.98 3.42 2.52 ;
        RECT  0.83 2.36 3.42 2.52 ;
        RECT  3.90 0.44 5.24 0.60 ;
        RECT  4.96 0.44 5.24 0.72 ;
        RECT  3.90 0.44 4.06 1.04 ;
        RECT  3.74 0.76 3.90 2.26 ;
        RECT  3.74 1.98 4.06 2.26 ;
        RECT  5.82 0.88 6.12 1.16 ;
        RECT  5.96 1.26 6.24 1.54 ;
        RECT  5.96 0.88 6.12 2.14 ;
        RECT  5.84 1.86 6.12 2.14 ;
        RECT  6.32 0.72 6.60 1.00 ;
        RECT  4.78 0.88 5.06 1.16 ;
        RECT  4.78 0.88 4.94 2.14 ;
        RECT  6.40 0.72 6.56 2.20 ;
        RECT  4.78 1.86 5.06 2.14 ;
        RECT  4.78 1.98 5.68 2.14 ;
        RECT  6.32 1.92 6.60 2.20 ;
        RECT  5.52 1.98 5.68 2.46 ;
        RECT  6.32 1.92 6.48 2.46 ;
        RECT  5.52 2.30 6.48 2.46 ;
        RECT  7.40 0.72 7.70 1.00 ;
        RECT  7.40 0.72 7.56 2.20 ;
        RECT  7.36 1.92 7.64 2.20 ;
        RECT  6.84 0.72 7.12 1.00 ;
        RECT  8.20 1.48 8.48 1.76 ;
        RECT  7.80 1.60 8.48 1.76 ;
        RECT  6.90 0.72 7.06 2.20 ;
        RECT  6.84 1.92 7.12 2.20 ;
        RECT  6.96 1.92 7.12 2.52 ;
        RECT  7.80 1.60 7.96 2.52 ;
        RECT  6.96 2.36 7.96 2.52 ;
        RECT  8.46 0.72 8.80 1.00 ;
        RECT  7.72 1.16 8.80 1.32 ;
        RECT  7.72 1.16 8.00 1.44 ;
        RECT  8.64 0.72 8.80 2.20 ;
        RECT  8.64 1.92 8.92 2.20 ;
        RECT  9.54 0.76 9.96 1.04 ;
        RECT  9.68 1.92 9.96 2.20 ;
        RECT  9.80 0.76 9.96 2.76 ;
        RECT  9.80 2.48 10.08 2.76 ;
        RECT  9.14 0.44 10.62 0.60 ;
        RECT  10.34 0.44 10.62 0.80 ;
        RECT  9.02 0.76 9.30 1.04 ;
        RECT  9.14 0.44 9.30 2.20 ;
        RECT  9.14 1.92 9.44 2.20 ;
        RECT  10.16 0.96 10.44 1.24 ;
        RECT  10.16 1.46 11.10 1.62 ;
        RECT  10.82 1.40 11.10 1.68 ;
        RECT  10.16 0.96 10.32 2.12 ;
        RECT  10.16 1.84 10.44 2.12 ;
        RECT  11.20 0.96 11.48 1.24 ;
        RECT  11.20 1.84 11.48 2.12 ;
        RECT  11.29 0.96 11.45 2.76 ;
        RECT  11.23 2.48 11.51 2.76 ;
    END
END DFFDEZSP4V1_0

MACRO DFFDEZSP2V1_0
    CLASS CORE ;
    FOREIGN DFFDEZSP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 13.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 25.20  LAYER ME1  ;
        ANTENNADIFFAREA 10.84  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.89  LAYER ME1  ;
        ANTENNAMAXAREACAR 28.22  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.72 1.90 13.00 2.18 ;
        RECT  12.72 0.96 13.00 1.24 ;
        RECT  12.72 0.96 12.88 2.18 ;
        RECT  12.46 1.46 12.88 1.74 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 25.20  LAYER ME1  ;
        ANTENNADIFFAREA 10.96  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.89  LAYER ME1  ;
        ANTENNAMAXAREACAR 28.22  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.21 1.88 1.51 2.16 ;
        RECT  1.21 0.66 1.51 0.96 ;
        RECT  1.21 0.66 1.37 2.16 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.99 1.46 2.34 1.76 ;
        END
    END E
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.45 1.06 2.78 1.34 ;
        RECT  2.26 1.06 2.78 1.30 ;
        END
    END SEL
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 25.20  LAYER ME1  ;
        ANTENNADIFFAREA 10.84  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.89  LAYER ME1  ;
        ANTENNAMAXAREACAR 28.22  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.68 1.90 11.96 2.18 ;
        RECT  11.68 0.96 11.96 1.24 ;
        RECT  11.69 0.96 11.94 2.18 ;
        RECT  11.66 1.46 11.94 1.74 ;
        END
    END Q
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.26 1.46 5.72 1.74 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 25.20  LAYER ME1  ;
        ANTENNADIFFAREA 10.96  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.89  LAYER ME1  ;
        ANTENNAMAXAREACAR 28.22  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.30 1.98 4.58 2.26 ;
        RECT  4.30 0.76 4.58 1.04 ;
        RECT  4.30 0.76 4.46 2.26 ;
        RECT  4.06 1.46 4.46 1.74 ;
        END
    END TD
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 13.20 0.28 ;
        RECT  12.74 -0.28 13.02 0.32 ;
        RECT  12.20 0.64 12.48 0.92 ;
        RECT  12.26 -0.28 12.42 0.92 ;
        RECT  10.68 0.96 10.96 1.24 ;
        RECT  10.78 -0.28 10.94 1.24 ;
        RECT  7.94 0.72 8.22 1.00 ;
        RECT  8.00 -0.28 8.16 1.00 ;
        RECT  5.30 0.88 5.58 1.16 ;
        RECT  5.40 -0.28 5.56 1.16 ;
        RECT  2.26 0.62 2.54 0.90 ;
        RECT  2.32 -0.28 2.48 0.90 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 13.20 3.48 ;
        RECT  12.74 2.88 13.02 3.48 ;
        RECT  12.20 2.22 12.48 2.50 ;
        RECT  12.26 2.22 12.42 3.48 ;
        RECT  10.68 1.84 10.96 2.12 ;
        RECT  10.74 1.84 10.90 3.48 ;
        RECT  8.12 1.92 8.40 2.20 ;
        RECT  8.18 1.92 8.34 3.48 ;
        RECT  5.09 2.52 5.37 3.48 ;
        RECT  3.78 2.52 4.06 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.19 0.68 0.47 0.96 ;
        RECT  0.19 1.88 0.47 2.16 ;
        RECT  0.19 0.68 0.35 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  1.67 0.62 2.02 0.90 ;
        RECT  1.53 1.12 1.83 1.40 ;
        RECT  1.67 0.62 1.83 2.20 ;
        RECT  1.67 1.92 2.02 2.20 ;
        RECT  2.78 0.62 3.10 0.90 ;
        RECT  2.94 1.22 3.22 1.50 ;
        RECT  2.94 0.62 3.10 2.20 ;
        RECT  2.78 1.92 3.10 2.20 ;
        RECT  0.71 0.68 0.99 0.96 ;
        RECT  3.26 0.76 3.54 1.04 ;
        RECT  0.77 0.68 0.93 2.16 ;
        RECT  0.71 1.88 0.99 2.16 ;
        RECT  3.38 0.76 3.54 2.26 ;
        RECT  0.83 1.88 0.99 2.52 ;
        RECT  3.26 1.98 3.42 2.52 ;
        RECT  0.83 2.36 3.42 2.52 ;
        RECT  3.90 0.44 5.24 0.60 ;
        RECT  4.96 0.44 5.24 0.72 ;
        RECT  3.90 0.44 4.06 1.04 ;
        RECT  3.74 0.76 3.90 2.26 ;
        RECT  3.74 1.98 4.06 2.26 ;
        RECT  5.82 0.88 6.12 1.16 ;
        RECT  5.96 1.26 6.24 1.54 ;
        RECT  5.96 0.88 6.12 2.14 ;
        RECT  5.84 1.86 6.12 2.14 ;
        RECT  6.32 0.72 6.60 1.00 ;
        RECT  4.78 0.88 5.06 1.16 ;
        RECT  4.78 0.88 4.94 2.14 ;
        RECT  6.40 0.72 6.56 2.20 ;
        RECT  4.78 1.86 5.06 2.14 ;
        RECT  4.78 1.98 5.68 2.14 ;
        RECT  6.32 1.92 6.60 2.20 ;
        RECT  5.52 1.98 5.68 2.46 ;
        RECT  6.32 1.92 6.48 2.46 ;
        RECT  5.52 2.30 6.48 2.46 ;
        RECT  7.40 0.72 7.70 1.00 ;
        RECT  7.40 0.72 7.56 2.20 ;
        RECT  7.36 1.92 7.64 2.20 ;
        RECT  6.84 0.72 7.12 1.00 ;
        RECT  8.20 1.48 8.48 1.76 ;
        RECT  7.80 1.60 8.48 1.76 ;
        RECT  6.90 0.72 7.06 2.20 ;
        RECT  6.84 1.92 7.12 2.20 ;
        RECT  6.96 1.92 7.12 2.52 ;
        RECT  7.80 1.60 7.96 2.52 ;
        RECT  6.96 2.36 7.96 2.52 ;
        RECT  8.46 0.72 8.80 1.00 ;
        RECT  7.72 1.16 8.80 1.32 ;
        RECT  7.72 1.16 8.00 1.44 ;
        RECT  8.64 0.72 8.80 2.20 ;
        RECT  8.64 1.92 8.92 2.20 ;
        RECT  9.54 0.76 9.96 1.04 ;
        RECT  9.68 1.92 9.96 2.20 ;
        RECT  9.80 0.76 9.96 2.76 ;
        RECT  9.80 2.48 10.08 2.76 ;
        RECT  9.14 0.44 10.62 0.60 ;
        RECT  10.34 0.44 10.62 0.80 ;
        RECT  9.02 0.76 9.30 1.04 ;
        RECT  9.14 0.44 9.30 2.20 ;
        RECT  9.14 1.92 9.44 2.20 ;
        RECT  10.16 0.96 10.44 1.24 ;
        RECT  10.16 1.46 11.10 1.62 ;
        RECT  10.82 1.40 11.10 1.68 ;
        RECT  10.16 0.96 10.32 2.12 ;
        RECT  10.16 1.84 10.44 2.12 ;
        RECT  11.20 0.96 11.48 1.24 ;
        RECT  11.20 1.84 11.48 2.12 ;
        RECT  11.29 0.96 11.45 2.76 ;
        RECT  11.23 2.48 11.51 2.76 ;
    END
END DFFDEZSP2V1_0

MACRO DFFDEZSP1V1_0
    CLASS CORE ;
    FOREIGN DFFDEZSP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 13.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 25.30  LAYER ME1  ;
        ANTENNADIFFAREA 10.26  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.74  LAYER ME1  ;
        ANTENNAMAXAREACAR 34.23  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.21 1.88 1.51 2.16 ;
        RECT  1.21 0.66 1.51 0.96 ;
        RECT  1.21 0.66 1.37 2.16 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.26 1.46 5.72 1.74 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 25.30  LAYER ME1  ;
        ANTENNADIFFAREA 10.15  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.74  LAYER ME1  ;
        ANTENNAMAXAREACAR 34.23  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.72 1.90 13.00 2.18 ;
        RECT  12.72 0.96 13.00 1.24 ;
        RECT  12.72 0.96 12.88 2.18 ;
        RECT  12.46 1.46 12.88 1.74 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 25.30  LAYER ME1  ;
        ANTENNADIFFAREA 10.15  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.74  LAYER ME1  ;
        ANTENNAMAXAREACAR 34.23  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.68 1.90 11.96 2.18 ;
        RECT  11.68 0.96 11.96 1.24 ;
        RECT  11.69 0.96 11.94 2.18 ;
        RECT  11.66 1.46 11.94 1.74 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.99 1.46 2.34 1.76 ;
        END
    END E
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.45 1.06 2.78 1.34 ;
        RECT  2.26 1.06 2.78 1.30 ;
        END
    END SEL
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 25.30  LAYER ME1  ;
        ANTENNADIFFAREA 10.26  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.74  LAYER ME1  ;
        ANTENNAMAXAREACAR 34.23  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.30 1.98 4.58 2.26 ;
        RECT  4.30 0.76 4.58 1.04 ;
        RECT  4.30 0.76 4.46 2.26 ;
        RECT  4.06 1.46 4.46 1.74 ;
        END
    END TD
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 13.20 3.48 ;
        RECT  12.74 2.88 13.02 3.48 ;
        RECT  12.20 1.90 12.48 2.18 ;
        RECT  12.26 1.90 12.42 3.48 ;
        RECT  10.68 1.84 10.96 2.12 ;
        RECT  10.74 1.84 10.90 3.48 ;
        RECT  8.12 1.92 8.40 2.20 ;
        RECT  8.18 1.92 8.34 3.48 ;
        RECT  5.09 2.52 5.37 3.48 ;
        RECT  3.78 2.52 4.06 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 13.20 0.28 ;
        RECT  12.74 -0.28 13.02 0.32 ;
        RECT  12.20 0.96 12.48 1.24 ;
        RECT  12.26 -0.28 12.42 1.24 ;
        RECT  10.68 0.96 10.96 1.24 ;
        RECT  10.78 -0.28 10.94 1.24 ;
        RECT  7.94 0.72 8.22 1.00 ;
        RECT  8.00 -0.28 8.16 1.00 ;
        RECT  5.30 0.88 5.58 1.16 ;
        RECT  5.40 -0.28 5.56 1.16 ;
        RECT  2.26 0.62 2.54 0.90 ;
        RECT  2.32 -0.28 2.48 0.90 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.19 0.68 0.47 0.96 ;
        RECT  0.19 1.88 0.47 2.16 ;
        RECT  0.19 0.68 0.35 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  1.67 0.62 2.02 0.90 ;
        RECT  1.53 1.12 1.83 1.40 ;
        RECT  1.67 0.62 1.83 2.20 ;
        RECT  1.67 1.92 2.02 2.20 ;
        RECT  2.78 0.62 3.10 0.90 ;
        RECT  2.94 1.22 3.22 1.50 ;
        RECT  2.94 0.62 3.10 2.20 ;
        RECT  2.78 1.92 3.10 2.20 ;
        RECT  0.71 0.68 0.99 0.96 ;
        RECT  3.26 0.76 3.54 1.04 ;
        RECT  0.77 0.68 0.93 2.16 ;
        RECT  0.71 1.88 0.99 2.16 ;
        RECT  3.38 0.76 3.54 2.26 ;
        RECT  0.83 1.88 0.99 2.52 ;
        RECT  3.26 1.98 3.42 2.52 ;
        RECT  0.83 2.36 3.42 2.52 ;
        RECT  3.90 0.44 5.24 0.60 ;
        RECT  4.96 0.44 5.24 0.72 ;
        RECT  3.90 0.44 4.06 1.04 ;
        RECT  3.74 0.76 3.90 2.26 ;
        RECT  3.74 1.98 4.06 2.26 ;
        RECT  5.82 0.88 6.12 1.16 ;
        RECT  5.96 1.26 6.24 1.54 ;
        RECT  5.96 0.88 6.12 2.14 ;
        RECT  5.84 1.86 6.12 2.14 ;
        RECT  6.32 0.72 6.60 1.00 ;
        RECT  4.78 0.88 5.06 1.16 ;
        RECT  4.78 0.88 4.94 2.14 ;
        RECT  6.40 0.72 6.56 2.20 ;
        RECT  4.78 1.86 5.06 2.14 ;
        RECT  4.78 1.98 5.68 2.14 ;
        RECT  6.32 1.92 6.60 2.20 ;
        RECT  5.52 1.98 5.68 2.46 ;
        RECT  6.32 1.92 6.48 2.46 ;
        RECT  5.52 2.30 6.48 2.46 ;
        RECT  7.40 0.72 7.70 1.00 ;
        RECT  7.40 0.72 7.56 2.20 ;
        RECT  7.36 1.92 7.64 2.20 ;
        RECT  6.84 0.72 7.12 1.00 ;
        RECT  8.20 1.48 8.48 1.76 ;
        RECT  7.80 1.60 8.48 1.76 ;
        RECT  6.90 0.72 7.06 2.20 ;
        RECT  6.84 1.92 7.12 2.20 ;
        RECT  6.96 1.92 7.12 2.52 ;
        RECT  7.80 1.60 7.96 2.52 ;
        RECT  6.96 2.36 7.96 2.52 ;
        RECT  8.46 0.72 8.80 1.00 ;
        RECT  7.72 1.16 8.80 1.32 ;
        RECT  7.72 1.16 8.00 1.44 ;
        RECT  8.64 0.72 8.80 2.20 ;
        RECT  8.64 1.92 8.92 2.20 ;
        RECT  9.54 0.76 9.96 1.04 ;
        RECT  9.68 1.92 9.96 2.20 ;
        RECT  9.80 0.76 9.96 2.76 ;
        RECT  9.80 2.48 10.08 2.76 ;
        RECT  9.14 0.44 10.62 0.60 ;
        RECT  10.34 0.44 10.62 0.80 ;
        RECT  9.02 0.76 9.30 1.04 ;
        RECT  9.14 0.44 9.30 2.20 ;
        RECT  9.14 1.92 9.44 2.20 ;
        RECT  10.16 0.96 10.44 1.24 ;
        RECT  10.16 1.46 11.10 1.62 ;
        RECT  10.82 1.40 11.10 1.68 ;
        RECT  10.16 0.96 10.32 2.12 ;
        RECT  10.16 1.84 10.44 2.12 ;
        RECT  11.20 0.96 11.48 1.24 ;
        RECT  11.20 1.84 11.48 2.12 ;
        RECT  11.29 0.96 11.45 2.76 ;
        RECT  11.23 2.48 11.51 2.76 ;
    END
END DFFDEZSP1V1_0

MACRO DFFDESZSP8V1_0
    CLASS CORE ;
    FOREIGN DFFDESZSP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 37.02  LAYER ME1  ;
        ANTENNADIFFAREA 17.59  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.76  LAYER ME1  ;
        ANTENNAMAXAREACAR 21.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  17.60 1.90 17.88 2.50 ;
        RECT  17.60 0.64 17.88 1.24 ;
        RECT  17.60 0.64 17.76 2.50 ;
        RECT  16.68 1.52 17.76 1.68 ;
        RECT  16.68 1.46 17.14 1.74 ;
        RECT  16.56 1.90 16.84 2.50 ;
        RECT  16.68 0.64 16.84 2.50 ;
        RECT  16.56 0.64 16.84 1.24 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 37.02  LAYER ME1  ;
        ANTENNADIFFAREA 17.56  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.76  LAYER ME1  ;
        ANTENNAMAXAREACAR 21.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  15.52 1.90 15.80 2.50 ;
        RECT  15.52 0.64 15.80 1.24 ;
        RECT  15.52 0.64 15.68 2.50 ;
        RECT  14.46 1.52 15.68 1.68 ;
        RECT  14.48 1.90 14.76 2.50 ;
        RECT  14.48 0.64 14.76 1.24 ;
        RECT  14.48 0.64 14.74 2.50 ;
        RECT  14.46 1.46 14.74 1.74 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 36.70  LAYER ME1  ;
        ANTENNADIFFAREA 16.98  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.76  LAYER ME1  ;
        ANTENNAMAXAREACAR 20.89  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.21 1.88 1.51 2.16 ;
        RECT  1.21 0.66 1.51 0.96 ;
        RECT  1.21 0.66 1.37 2.16 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.99 1.46 2.34 1.76 ;
        END
    END E
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.92 1.40 12.34 1.68 ;
        END
    END SB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.64 1.40 5.94 1.76 ;
        END
    END CK
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.45 1.06 2.78 1.34 ;
        RECT  2.26 1.06 2.78 1.30 ;
        END
    END SEL
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 37.02  LAYER ME1  ;
        ANTENNADIFFAREA 16.98  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.76  LAYER ME1  ;
        ANTENNAMAXAREACAR 21.07  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.42 1.46 4.74 1.74 ;
        RECT  4.34 0.88 4.62 1.16 ;
        RECT  4.30 1.98 4.58 2.26 ;
        RECT  4.42 0.88 4.58 2.26 ;
        END
    END TD
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 18.80 0.28 ;
        RECT  18.18 -0.28 18.62 0.32 ;
        RECT  18.12 0.64 18.40 1.24 ;
        RECT  18.18 -0.28 18.34 1.24 ;
        RECT  17.08 0.64 17.36 1.24 ;
        RECT  17.14 -0.28 17.30 1.24 ;
        RECT  16.04 0.64 16.32 1.24 ;
        RECT  16.10 -0.28 16.26 1.24 ;
        RECT  15.00 0.64 15.28 1.24 ;
        RECT  15.06 -0.28 15.22 1.24 ;
        RECT  13.96 0.64 14.24 1.24 ;
        RECT  14.02 -0.28 14.18 1.24 ;
        RECT  12.96 0.88 13.24 1.16 ;
        RECT  13.02 -0.28 13.18 1.16 ;
        RECT  11.48 -0.28 11.76 0.68 ;
        RECT  5.06 -0.28 5.34 0.64 ;
        RECT  2.26 0.62 2.54 0.90 ;
        RECT  2.32 -0.28 2.48 0.90 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 18.80 3.48 ;
        RECT  18.18 2.88 18.62 3.48 ;
        RECT  18.12 1.90 18.40 2.50 ;
        RECT  18.18 1.90 18.34 3.48 ;
        RECT  17.08 1.90 17.36 2.50 ;
        RECT  17.14 1.90 17.30 3.48 ;
        RECT  16.04 1.90 16.32 2.50 ;
        RECT  16.10 1.90 16.26 3.48 ;
        RECT  15.00 1.90 15.28 2.50 ;
        RECT  15.06 1.90 15.22 3.48 ;
        RECT  13.96 1.90 14.24 2.50 ;
        RECT  14.02 1.90 14.18 3.48 ;
        RECT  12.72 2.40 13.00 3.48 ;
        RECT  11.92 1.84 12.20 2.12 ;
        RECT  11.98 1.84 12.14 3.48 ;
        RECT  10.92 1.84 11.20 2.12 ;
        RECT  10.98 1.84 11.14 3.48 ;
        RECT  9.92 1.84 10.20 2.12 ;
        RECT  10.02 1.84 10.18 3.48 ;
        RECT  5.06 2.52 5.34 3.48 ;
        RECT  3.78 2.52 4.06 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.19 0.68 0.47 0.96 ;
        RECT  0.19 1.88 0.47 2.16 ;
        RECT  0.19 0.68 0.35 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  1.67 0.62 2.02 0.90 ;
        RECT  1.53 1.12 1.83 1.40 ;
        RECT  1.67 0.62 1.83 2.20 ;
        RECT  1.67 1.92 2.02 2.20 ;
        RECT  2.78 0.62 3.10 0.90 ;
        RECT  2.94 1.22 3.22 1.50 ;
        RECT  2.94 0.62 3.10 2.20 ;
        RECT  2.78 1.92 3.10 2.20 ;
        RECT  0.71 0.68 0.99 0.96 ;
        RECT  3.26 0.76 3.54 1.04 ;
        RECT  0.77 0.68 0.93 2.16 ;
        RECT  0.71 1.88 0.99 2.16 ;
        RECT  3.38 0.76 3.54 2.26 ;
        RECT  0.83 1.88 0.99 2.52 ;
        RECT  3.26 1.98 3.42 2.52 ;
        RECT  0.83 2.36 3.42 2.52 ;
        RECT  3.90 0.44 4.90 0.60 ;
        RECT  4.62 0.44 4.90 0.72 ;
        RECT  3.90 0.44 4.06 1.04 ;
        RECT  3.74 0.76 3.90 2.26 ;
        RECT  3.74 1.98 4.06 2.26 ;
        RECT  5.82 0.96 6.26 1.24 ;
        RECT  6.10 1.46 6.42 1.74 ;
        RECT  6.10 0.96 6.26 2.20 ;
        RECT  5.82 1.92 6.26 2.20 ;
        RECT  6.42 0.44 6.70 0.72 ;
        RECT  5.50 0.56 6.70 0.72 ;
        RECT  5.50 0.56 5.66 1.12 ;
        RECT  4.82 0.96 5.66 1.12 ;
        RECT  4.82 0.96 5.10 1.24 ;
        RECT  4.90 0.96 5.06 2.20 ;
        RECT  4.78 1.92 5.06 2.20 ;
        RECT  4.78 2.04 5.66 2.20 ;
        RECT  5.50 2.04 5.66 2.64 ;
        RECT  5.50 2.48 6.60 2.64 ;
        RECT  6.32 2.48 6.60 2.76 ;
        RECT  7.94 0.76 8.26 1.04 ;
        RECT  7.94 0.76 8.10 2.00 ;
        RECT  7.60 1.84 8.64 2.00 ;
        RECT  7.60 1.84 7.88 2.12 ;
        RECT  8.36 1.84 8.64 2.12 ;
        RECT  8.50 0.76 8.78 1.04 ;
        RECT  8.62 0.76 8.78 1.36 ;
        RECT  9.46 1.08 9.74 1.36 ;
        RECT  8.62 1.20 9.74 1.36 ;
        RECT  8.88 1.20 9.04 2.12 ;
        RECT  8.88 1.84 9.16 2.12 ;
        RECT  6.98 0.86 7.26 1.14 ;
        RECT  6.42 0.98 7.26 1.14 ;
        RECT  6.42 0.96 6.70 1.24 ;
        RECT  6.64 0.98 6.80 2.12 ;
        RECT  6.76 1.84 6.92 2.44 ;
        RECT  6.76 2.28 9.86 2.44 ;
        RECT  9.58 2.28 9.86 2.56 ;
        RECT  9.02 0.76 10.30 0.92 ;
        RECT  9.02 0.76 9.30 1.04 ;
        RECT  10.02 0.76 10.30 1.16 ;
        RECT  10.02 0.76 10.18 1.68 ;
        RECT  11.06 1.40 11.34 1.68 ;
        RECT  9.60 1.52 11.34 1.68 ;
        RECT  10.36 1.52 10.52 2.12 ;
        RECT  9.60 1.52 9.76 2.12 ;
        RECT  9.40 1.84 9.76 2.12 ;
        RECT  10.36 1.84 10.72 2.12 ;
        RECT  7.62 0.44 11.22 0.60 ;
        RECT  11.06 0.44 11.22 1.04 ;
        RECT  11.06 0.88 11.72 1.04 ;
        RECT  7.62 0.44 7.78 1.14 ;
        RECT  11.44 0.88 11.72 1.16 ;
        RECT  7.50 0.86 7.66 1.46 ;
        RECT  7.28 1.30 7.66 1.46 ;
        RECT  11.50 0.88 11.66 2.12 ;
        RECT  7.28 1.30 7.44 2.12 ;
        RECT  7.16 1.84 7.44 2.12 ;
        RECT  11.44 1.84 11.72 2.12 ;
        RECT  12.06 0.88 12.34 1.16 ;
        RECT  12.06 1.00 12.66 1.16 ;
        RECT  12.50 1.00 12.66 2.12 ;
        RECT  12.44 1.84 12.72 2.12 ;
        RECT  12.44 1.96 13.32 2.12 ;
        RECT  13.16 1.96 13.32 2.64 ;
        RECT  13.16 2.48 13.79 2.64 ;
        RECT  13.51 2.48 13.79 2.76 ;
        RECT  13.48 0.88 13.76 1.16 ;
        RECT  12.82 1.46 13.90 1.62 ;
        RECT  12.82 1.40 13.10 1.68 ;
        RECT  13.60 1.40 13.90 1.68 ;
        RECT  13.60 0.88 13.76 2.12 ;
        RECT  13.48 1.84 13.76 2.12 ;
    END
END DFFDESZSP8V1_0

MACRO DFFDESZSP4V1_0
    CLASS CORE ;
    FOREIGN DFFDESZSP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.64 1.40 5.94 1.76 ;
        END
    END CK
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.92 1.40 12.34 1.68 ;
        END
    END SB
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.99 1.46 2.34 1.76 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 32.43  LAYER ME1  ;
        ANTENNADIFFAREA 14.42  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.18  LAYER ME1  ;
        ANTENNAMAXAREACAR 27.47  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.21 1.88 1.51 2.16 ;
        RECT  1.21 0.66 1.51 0.96 ;
        RECT  1.21 0.66 1.37 2.16 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 32.75  LAYER ME1  ;
        ANTENNADIFFAREA 14.52  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.18  LAYER ME1  ;
        ANTENNAMAXAREACAR 27.74  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.48 1.90 14.76 2.50 ;
        RECT  14.48 0.64 14.76 1.24 ;
        RECT  14.48 0.64 14.74 2.50 ;
        RECT  14.46 1.46 14.74 1.74 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 32.75  LAYER ME1  ;
        ANTENNADIFFAREA 14.55  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.18  LAYER ME1  ;
        ANTENNAMAXAREACAR 27.74  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  15.64 1.46 15.94 1.74 ;
        RECT  15.52 1.90 15.80 2.50 ;
        RECT  15.64 0.64 15.80 2.50 ;
        RECT  15.52 0.64 15.80 1.24 ;
        END
    END QB
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.45 1.06 2.78 1.34 ;
        RECT  2.26 1.06 2.78 1.30 ;
        END
    END SEL
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 32.75  LAYER ME1  ;
        ANTENNADIFFAREA 14.42  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.18  LAYER ME1  ;
        ANTENNAMAXAREACAR 27.74  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.42 1.46 4.74 1.74 ;
        RECT  4.34 0.88 4.62 1.16 ;
        RECT  4.30 1.98 4.58 2.26 ;
        RECT  4.42 0.88 4.58 2.26 ;
        END
    END TD
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 16.80 3.48 ;
        RECT  16.18 2.88 16.62 3.48 ;
        RECT  16.18 1.90 16.34 3.48 ;
        RECT  16.04 1.90 16.34 2.50 ;
        RECT  15.00 1.90 15.28 2.50 ;
        RECT  15.06 1.90 15.22 3.48 ;
        RECT  13.96 1.90 14.24 2.50 ;
        RECT  14.02 1.90 14.18 3.48 ;
        RECT  12.72 2.40 13.00 3.48 ;
        RECT  11.92 1.84 12.20 2.12 ;
        RECT  11.98 1.84 12.14 3.48 ;
        RECT  10.92 1.84 11.20 2.12 ;
        RECT  10.98 1.84 11.14 3.48 ;
        RECT  9.92 1.84 10.20 2.12 ;
        RECT  10.02 1.84 10.18 3.48 ;
        RECT  5.06 2.52 5.34 3.48 ;
        RECT  3.78 2.52 4.06 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 16.80 0.28 ;
        RECT  16.18 -0.28 16.62 0.32 ;
        RECT  16.04 0.64 16.34 1.24 ;
        RECT  16.18 -0.28 16.34 1.24 ;
        RECT  15.00 0.64 15.28 1.24 ;
        RECT  15.06 -0.28 15.22 1.24 ;
        RECT  13.96 0.64 14.24 1.24 ;
        RECT  14.02 -0.28 14.18 1.24 ;
        RECT  12.96 0.88 13.24 1.16 ;
        RECT  13.02 -0.28 13.18 1.16 ;
        RECT  11.48 -0.28 11.76 0.68 ;
        RECT  5.06 -0.28 5.34 0.64 ;
        RECT  2.26 0.62 2.54 0.90 ;
        RECT  2.32 -0.28 2.48 0.90 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.19 0.68 0.47 0.96 ;
        RECT  0.19 1.88 0.47 2.16 ;
        RECT  0.19 0.68 0.35 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  1.67 0.62 2.02 0.90 ;
        RECT  1.53 1.12 1.83 1.40 ;
        RECT  1.67 0.62 1.83 2.20 ;
        RECT  1.67 1.92 2.02 2.20 ;
        RECT  2.78 0.62 3.10 0.90 ;
        RECT  2.94 1.22 3.22 1.50 ;
        RECT  2.94 0.62 3.10 2.20 ;
        RECT  2.78 1.92 3.10 2.20 ;
        RECT  0.71 0.68 0.99 0.96 ;
        RECT  3.26 0.76 3.54 1.04 ;
        RECT  0.77 0.68 0.93 2.16 ;
        RECT  0.71 1.88 0.99 2.16 ;
        RECT  3.38 0.76 3.54 2.26 ;
        RECT  0.83 1.88 0.99 2.52 ;
        RECT  3.26 1.98 3.42 2.52 ;
        RECT  0.83 2.36 3.42 2.52 ;
        RECT  3.90 0.44 4.90 0.60 ;
        RECT  4.62 0.44 4.90 0.72 ;
        RECT  3.90 0.44 4.06 1.04 ;
        RECT  3.74 0.76 3.90 2.26 ;
        RECT  3.74 1.98 4.06 2.26 ;
        RECT  5.82 0.96 6.26 1.24 ;
        RECT  6.10 1.46 6.42 1.74 ;
        RECT  6.10 0.96 6.26 2.20 ;
        RECT  5.82 1.92 6.26 2.20 ;
        RECT  6.42 0.44 6.70 0.72 ;
        RECT  5.50 0.56 6.70 0.72 ;
        RECT  5.50 0.56 5.66 1.12 ;
        RECT  4.82 0.96 5.66 1.12 ;
        RECT  4.82 0.96 5.10 1.24 ;
        RECT  4.90 0.96 5.06 2.20 ;
        RECT  4.78 1.92 5.06 2.20 ;
        RECT  4.78 2.04 5.66 2.20 ;
        RECT  5.50 2.04 5.66 2.64 ;
        RECT  5.50 2.48 6.60 2.64 ;
        RECT  6.32 2.48 6.60 2.76 ;
        RECT  7.94 0.76 8.26 1.04 ;
        RECT  7.94 0.76 8.10 2.00 ;
        RECT  7.60 1.84 8.64 2.00 ;
        RECT  7.60 1.84 7.88 2.12 ;
        RECT  8.36 1.84 8.64 2.12 ;
        RECT  8.50 0.76 8.78 1.04 ;
        RECT  8.62 0.76 8.78 1.36 ;
        RECT  9.46 1.08 9.74 1.36 ;
        RECT  8.62 1.20 9.74 1.36 ;
        RECT  8.88 1.20 9.04 2.12 ;
        RECT  8.88 1.84 9.16 2.12 ;
        RECT  6.98 0.86 7.26 1.14 ;
        RECT  6.42 0.98 7.26 1.14 ;
        RECT  6.42 0.96 6.70 1.24 ;
        RECT  6.64 0.98 6.80 2.12 ;
        RECT  6.76 1.84 6.92 2.44 ;
        RECT  6.76 2.28 9.86 2.44 ;
        RECT  9.58 2.28 9.86 2.56 ;
        RECT  9.02 0.76 10.30 0.92 ;
        RECT  9.02 0.76 9.30 1.04 ;
        RECT  10.02 0.76 10.30 1.16 ;
        RECT  10.02 0.76 10.18 1.68 ;
        RECT  11.06 1.40 11.34 1.68 ;
        RECT  9.60 1.52 11.34 1.68 ;
        RECT  10.36 1.52 10.52 2.12 ;
        RECT  9.60 1.52 9.76 2.12 ;
        RECT  9.40 1.84 9.76 2.12 ;
        RECT  10.36 1.84 10.72 2.12 ;
        RECT  7.62 0.44 11.22 0.60 ;
        RECT  11.06 0.44 11.22 1.04 ;
        RECT  11.06 0.88 11.72 1.04 ;
        RECT  7.62 0.44 7.78 1.14 ;
        RECT  11.44 0.88 11.72 1.16 ;
        RECT  7.50 0.86 7.66 1.46 ;
        RECT  7.28 1.30 7.66 1.46 ;
        RECT  11.50 0.88 11.66 2.12 ;
        RECT  7.28 1.30 7.44 2.12 ;
        RECT  7.16 1.84 7.44 2.12 ;
        RECT  11.44 1.84 11.72 2.12 ;
        RECT  12.06 0.88 12.34 1.16 ;
        RECT  12.06 1.00 12.66 1.16 ;
        RECT  12.50 1.00 12.66 2.12 ;
        RECT  12.44 1.84 12.72 2.12 ;
        RECT  12.44 1.96 13.32 2.12 ;
        RECT  13.16 1.96 13.32 2.64 ;
        RECT  13.16 2.48 13.79 2.64 ;
        RECT  13.51 2.48 13.79 2.76 ;
        RECT  13.48 0.88 13.76 1.16 ;
        RECT  12.82 1.46 13.90 1.62 ;
        RECT  12.82 1.40 13.10 1.68 ;
        RECT  13.60 1.40 13.90 1.68 ;
        RECT  13.60 0.88 13.76 2.12 ;
        RECT  13.48 1.84 13.76 2.12 ;
    END
END DFFDESZSP4V1_0

MACRO DFFDESZSP2V1_0
    CLASS CORE ;
    FOREIGN DFFDESZSP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 30.46  LAYER ME1  ;
        ANTENNADIFFAREA 12.97  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.89  LAYER ME1  ;
        ANTENNAMAXAREACAR 34.12  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  15.12 1.46 15.52 1.74 ;
        RECT  15.00 1.90 15.28 2.50 ;
        RECT  15.12 0.64 15.28 2.50 ;
        RECT  15.00 0.64 15.28 1.24 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 30.46  LAYER ME1  ;
        ANTENNADIFFAREA 12.97  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.89  LAYER ME1  ;
        ANTENNAMAXAREACAR 34.12  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.06 1.46 14.34 1.74 ;
        RECT  13.96 1.90 14.24 2.50 ;
        RECT  14.06 0.64 14.24 2.50 ;
        RECT  13.96 0.64 14.24 1.24 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 30.14  LAYER ME1  ;
        ANTENNADIFFAREA 13.08  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.89  LAYER ME1  ;
        ANTENNAMAXAREACAR 33.76  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.21 1.88 1.51 2.16 ;
        RECT  1.21 0.66 1.51 0.96 ;
        RECT  1.21 0.66 1.37 2.16 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.99 1.46 2.34 1.76 ;
        END
    END E
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.92 1.40 12.34 1.68 ;
        END
    END SB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.64 1.40 5.94 1.76 ;
        END
    END CK
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.45 1.06 2.78 1.34 ;
        RECT  2.26 1.06 2.78 1.30 ;
        END
    END SEL
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 30.46  LAYER ME1  ;
        ANTENNADIFFAREA 13.08  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.89  LAYER ME1  ;
        ANTENNAMAXAREACAR 34.12  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.42 1.46 4.74 1.74 ;
        RECT  4.34 0.88 4.62 1.16 ;
        RECT  4.30 1.98 4.58 2.26 ;
        RECT  4.42 0.88 4.58 2.26 ;
        END
    END TD
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 15.60 0.28 ;
        RECT  15.14 -0.28 15.42 0.32 ;
        RECT  14.48 0.64 14.76 1.24 ;
        RECT  14.54 -0.28 14.70 1.24 ;
        RECT  12.96 0.88 13.24 1.16 ;
        RECT  13.02 -0.28 13.18 1.16 ;
        RECT  11.48 -0.28 11.76 0.68 ;
        RECT  5.06 -0.28 5.34 0.64 ;
        RECT  2.26 0.62 2.54 0.90 ;
        RECT  2.32 -0.28 2.48 0.90 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 15.60 3.48 ;
        RECT  15.14 2.88 15.42 3.48 ;
        RECT  14.48 1.90 14.76 2.50 ;
        RECT  14.54 1.90 14.70 3.48 ;
        RECT  12.72 2.40 13.00 3.48 ;
        RECT  11.92 1.84 12.20 2.12 ;
        RECT  11.98 1.84 12.14 3.48 ;
        RECT  10.92 1.84 11.20 2.12 ;
        RECT  10.98 1.84 11.14 3.48 ;
        RECT  9.92 1.84 10.20 2.12 ;
        RECT  10.02 1.84 10.18 3.48 ;
        RECT  5.06 2.52 5.34 3.48 ;
        RECT  3.78 2.52 4.06 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.19 0.68 0.47 0.96 ;
        RECT  0.19 1.88 0.47 2.16 ;
        RECT  0.19 0.68 0.35 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  1.67 0.62 2.02 0.90 ;
        RECT  1.53 1.12 1.83 1.40 ;
        RECT  1.67 0.62 1.83 2.20 ;
        RECT  1.67 1.92 2.02 2.20 ;
        RECT  2.78 0.62 3.10 0.90 ;
        RECT  2.94 1.22 3.22 1.50 ;
        RECT  2.94 0.62 3.10 2.20 ;
        RECT  2.78 1.92 3.10 2.20 ;
        RECT  0.71 0.68 0.99 0.96 ;
        RECT  3.26 0.76 3.54 1.04 ;
        RECT  0.77 0.68 0.93 2.16 ;
        RECT  0.71 1.88 0.99 2.16 ;
        RECT  3.38 0.76 3.54 2.26 ;
        RECT  0.83 1.88 0.99 2.52 ;
        RECT  3.26 1.98 3.42 2.52 ;
        RECT  0.83 2.36 3.42 2.52 ;
        RECT  3.90 0.44 4.90 0.60 ;
        RECT  4.62 0.44 4.90 0.72 ;
        RECT  3.90 0.44 4.06 1.04 ;
        RECT  3.74 0.76 3.90 2.26 ;
        RECT  3.74 1.98 4.06 2.26 ;
        RECT  5.82 0.96 6.26 1.24 ;
        RECT  6.10 1.46 6.42 1.74 ;
        RECT  6.10 0.96 6.26 2.20 ;
        RECT  5.82 1.92 6.26 2.20 ;
        RECT  6.42 0.44 6.70 0.72 ;
        RECT  5.50 0.56 6.70 0.72 ;
        RECT  5.50 0.56 5.66 1.12 ;
        RECT  4.82 0.96 5.66 1.12 ;
        RECT  4.82 0.96 5.10 1.24 ;
        RECT  4.90 0.96 5.06 2.20 ;
        RECT  4.78 1.92 5.06 2.20 ;
        RECT  4.78 2.04 5.66 2.20 ;
        RECT  5.50 2.04 5.66 2.64 ;
        RECT  5.50 2.48 6.60 2.64 ;
        RECT  6.32 2.48 6.60 2.76 ;
        RECT  7.94 0.76 8.26 1.04 ;
        RECT  7.94 0.76 8.10 2.00 ;
        RECT  7.60 1.84 8.64 2.00 ;
        RECT  7.60 1.84 7.88 2.12 ;
        RECT  8.36 1.84 8.64 2.12 ;
        RECT  8.50 0.76 8.78 1.04 ;
        RECT  8.62 0.76 8.78 1.36 ;
        RECT  9.46 1.08 9.74 1.36 ;
        RECT  8.62 1.20 9.74 1.36 ;
        RECT  8.88 1.20 9.04 2.12 ;
        RECT  8.88 1.84 9.16 2.12 ;
        RECT  6.98 0.86 7.26 1.14 ;
        RECT  6.42 0.98 7.26 1.14 ;
        RECT  6.42 0.96 6.70 1.24 ;
        RECT  6.64 0.98 6.80 2.12 ;
        RECT  6.76 1.84 6.92 2.44 ;
        RECT  6.76 2.28 9.86 2.44 ;
        RECT  9.58 2.28 9.86 2.56 ;
        RECT  9.02 0.76 10.30 0.92 ;
        RECT  9.02 0.76 9.30 1.04 ;
        RECT  10.02 0.76 10.30 1.16 ;
        RECT  10.02 0.76 10.18 1.68 ;
        RECT  11.06 1.40 11.34 1.68 ;
        RECT  9.60 1.52 11.34 1.68 ;
        RECT  10.36 1.52 10.52 2.12 ;
        RECT  9.60 1.52 9.76 2.12 ;
        RECT  9.40 1.84 9.76 2.12 ;
        RECT  10.36 1.84 10.72 2.12 ;
        RECT  7.62 0.44 11.22 0.60 ;
        RECT  11.06 0.44 11.22 1.04 ;
        RECT  11.06 0.88 11.72 1.04 ;
        RECT  7.62 0.44 7.78 1.14 ;
        RECT  11.44 0.88 11.72 1.16 ;
        RECT  7.50 0.86 7.66 1.46 ;
        RECT  7.28 1.30 7.66 1.46 ;
        RECT  11.50 0.88 11.66 2.12 ;
        RECT  7.28 1.30 7.44 2.12 ;
        RECT  7.16 1.84 7.44 2.12 ;
        RECT  11.44 1.84 11.72 2.12 ;
        RECT  12.06 0.88 12.34 1.16 ;
        RECT  12.06 1.00 12.66 1.16 ;
        RECT  12.50 1.00 12.66 2.12 ;
        RECT  12.44 1.84 12.72 2.12 ;
        RECT  12.44 1.96 13.32 2.12 ;
        RECT  13.16 1.96 13.32 2.64 ;
        RECT  13.16 2.48 13.79 2.64 ;
        RECT  13.51 2.48 13.79 2.76 ;
        RECT  13.48 0.88 13.76 1.16 ;
        RECT  12.82 1.46 13.90 1.62 ;
        RECT  12.82 1.40 13.10 1.68 ;
        RECT  13.60 1.40 13.90 1.68 ;
        RECT  13.60 0.88 13.76 2.12 ;
        RECT  13.48 1.84 13.76 2.12 ;
    END
END DFFDESZSP2V1_0

MACRO DFFDESZSP1V1_0
    CLASS CORE ;
    FOREIGN DFFDESZSP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.64 1.40 5.94 1.76 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 30.03  LAYER ME1  ;
        ANTENNADIFFAREA 12.28  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.74  LAYER ME1  ;
        ANTENNAMAXAREACAR 40.62  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  15.12 1.46 15.52 1.74 ;
        RECT  15.00 1.90 15.28 2.18 ;
        RECT  15.12 0.96 15.28 2.18 ;
        RECT  15.00 0.96 15.28 1.24 ;
        END
    END QB
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.92 1.40 12.34 1.68 ;
        END
    END SB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 29.72  LAYER ME1  ;
        ANTENNADIFFAREA 12.28  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.74  LAYER ME1  ;
        ANTENNAMAXAREACAR 40.21  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.06 1.46 14.34 1.74 ;
        RECT  13.96 1.90 14.24 2.18 ;
        RECT  14.06 0.96 14.24 2.18 ;
        RECT  13.96 0.96 14.24 1.24 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.99 1.46 2.34 1.76 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 30.03  LAYER ME1  ;
        ANTENNADIFFAREA 12.39  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.74  LAYER ME1  ;
        ANTENNAMAXAREACAR 40.62  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.21 1.88 1.51 2.16 ;
        RECT  1.21 0.66 1.51 0.96 ;
        RECT  1.21 0.66 1.37 2.16 ;
        END
    END D
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 30.03  LAYER ME1  ;
        ANTENNADIFFAREA 12.39  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.74  LAYER ME1  ;
        ANTENNAMAXAREACAR 40.62  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.42 1.46 4.74 1.74 ;
        RECT  4.34 0.88 4.62 1.16 ;
        RECT  4.30 1.98 4.58 2.26 ;
        RECT  4.42 0.88 4.58 2.26 ;
        END
    END TD
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.45 1.06 2.78 1.34 ;
        RECT  2.26 1.06 2.78 1.30 ;
        END
    END SEL
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 15.60 0.28 ;
        RECT  15.14 -0.28 15.42 0.32 ;
        RECT  14.48 0.96 14.76 1.24 ;
        RECT  14.54 -0.28 14.70 1.24 ;
        RECT  12.96 0.88 13.24 1.16 ;
        RECT  13.02 -0.28 13.18 1.16 ;
        RECT  11.48 -0.28 11.76 0.68 ;
        RECT  5.06 -0.28 5.34 0.64 ;
        RECT  2.26 0.62 2.54 0.90 ;
        RECT  2.32 -0.28 2.48 0.90 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 15.60 3.48 ;
        RECT  15.14 2.88 15.42 3.48 ;
        RECT  14.48 1.90 14.76 2.18 ;
        RECT  14.54 1.90 14.70 3.48 ;
        RECT  12.72 2.40 13.00 3.48 ;
        RECT  11.92 1.84 12.20 2.12 ;
        RECT  11.98 1.84 12.14 3.48 ;
        RECT  10.92 1.84 11.20 2.12 ;
        RECT  10.98 1.84 11.14 3.48 ;
        RECT  9.92 1.84 10.20 2.12 ;
        RECT  10.02 1.84 10.18 3.48 ;
        RECT  5.06 2.52 5.34 3.48 ;
        RECT  3.78 2.52 4.06 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.19 0.68 0.47 0.96 ;
        RECT  0.19 1.88 0.47 2.16 ;
        RECT  0.19 0.68 0.35 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  1.67 0.62 2.02 0.90 ;
        RECT  1.53 1.12 1.83 1.40 ;
        RECT  1.67 0.62 1.83 2.20 ;
        RECT  1.67 1.92 2.02 2.20 ;
        RECT  2.78 0.62 3.10 0.90 ;
        RECT  2.94 1.22 3.22 1.50 ;
        RECT  2.94 0.62 3.10 2.20 ;
        RECT  2.78 1.92 3.10 2.20 ;
        RECT  0.71 0.68 0.99 0.96 ;
        RECT  3.26 0.76 3.54 1.04 ;
        RECT  0.77 0.68 0.93 2.16 ;
        RECT  0.71 1.88 0.99 2.16 ;
        RECT  3.38 0.76 3.54 2.26 ;
        RECT  0.83 1.88 0.99 2.52 ;
        RECT  3.26 1.98 3.42 2.52 ;
        RECT  0.83 2.36 3.42 2.52 ;
        RECT  3.90 0.44 4.90 0.60 ;
        RECT  4.62 0.44 4.90 0.72 ;
        RECT  3.90 0.44 4.06 1.04 ;
        RECT  3.74 0.76 3.90 2.26 ;
        RECT  3.74 1.98 4.06 2.26 ;
        RECT  5.82 0.96 6.26 1.24 ;
        RECT  6.10 1.46 6.42 1.74 ;
        RECT  6.10 0.96 6.26 2.20 ;
        RECT  5.82 1.92 6.26 2.20 ;
        RECT  6.42 0.44 6.70 0.72 ;
        RECT  5.50 0.56 6.70 0.72 ;
        RECT  5.50 0.56 5.66 1.12 ;
        RECT  4.82 0.96 5.66 1.12 ;
        RECT  4.82 0.96 5.10 1.24 ;
        RECT  4.90 0.96 5.06 2.20 ;
        RECT  4.78 1.92 5.06 2.20 ;
        RECT  4.78 2.04 5.66 2.20 ;
        RECT  5.50 2.04 5.66 2.64 ;
        RECT  5.50 2.48 6.60 2.64 ;
        RECT  6.32 2.48 6.60 2.76 ;
        RECT  7.94 0.76 8.26 1.04 ;
        RECT  7.94 0.76 8.10 2.00 ;
        RECT  7.60 1.84 8.64 2.00 ;
        RECT  7.60 1.84 7.88 2.12 ;
        RECT  8.36 1.84 8.64 2.12 ;
        RECT  8.50 0.76 8.78 1.04 ;
        RECT  8.62 0.76 8.78 1.36 ;
        RECT  9.46 1.08 9.74 1.36 ;
        RECT  8.62 1.20 9.74 1.36 ;
        RECT  8.88 1.20 9.04 2.12 ;
        RECT  8.88 1.84 9.16 2.12 ;
        RECT  6.98 0.86 7.26 1.14 ;
        RECT  6.42 0.98 7.26 1.14 ;
        RECT  6.42 0.96 6.70 1.24 ;
        RECT  6.64 0.98 6.80 2.12 ;
        RECT  6.76 1.84 6.92 2.44 ;
        RECT  6.76 2.28 9.86 2.44 ;
        RECT  9.58 2.28 9.86 2.56 ;
        RECT  9.02 0.76 10.30 0.92 ;
        RECT  9.02 0.76 9.30 1.04 ;
        RECT  10.02 0.76 10.30 1.16 ;
        RECT  10.02 0.76 10.18 1.68 ;
        RECT  11.06 1.40 11.34 1.68 ;
        RECT  9.60 1.52 11.34 1.68 ;
        RECT  10.36 1.52 10.52 2.12 ;
        RECT  9.60 1.52 9.76 2.12 ;
        RECT  9.40 1.84 9.76 2.12 ;
        RECT  10.36 1.84 10.72 2.12 ;
        RECT  7.62 0.44 11.22 0.60 ;
        RECT  11.06 0.44 11.22 1.04 ;
        RECT  11.06 0.88 11.72 1.04 ;
        RECT  7.62 0.44 7.78 1.14 ;
        RECT  11.44 0.88 11.72 1.16 ;
        RECT  7.50 0.86 7.66 1.46 ;
        RECT  7.28 1.30 7.66 1.46 ;
        RECT  11.50 0.88 11.66 2.12 ;
        RECT  7.28 1.30 7.44 2.12 ;
        RECT  7.16 1.84 7.44 2.12 ;
        RECT  11.44 1.84 11.72 2.12 ;
        RECT  12.06 0.88 12.34 1.16 ;
        RECT  12.06 1.00 12.66 1.16 ;
        RECT  12.50 1.00 12.66 2.12 ;
        RECT  12.44 1.84 12.72 2.12 ;
        RECT  12.44 1.96 13.32 2.12 ;
        RECT  13.16 1.96 13.32 2.64 ;
        RECT  13.16 2.48 13.79 2.64 ;
        RECT  13.51 2.48 13.79 2.76 ;
        RECT  13.48 0.88 13.76 1.16 ;
        RECT  12.82 1.46 13.90 1.62 ;
        RECT  12.82 1.40 13.10 1.68 ;
        RECT  13.60 1.40 13.90 1.68 ;
        RECT  13.60 0.88 13.76 2.12 ;
        RECT  13.48 1.84 13.76 2.12 ;
    END
END DFFDESZSP1V1_0

MACRO DFFDESSP8V1_0
    CLASS CORE ;
    FOREIGN DFFDESSP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.24 1.40 3.54 1.76 ;
        END
    END CK
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.53 1.40 9.95 1.68 ;
        END
    END SB
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 32.42  LAYER ME1  ;
        ANTENNADIFFAREA 15.01  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.69  LAYER ME1  ;
        ANTENNAMAXAREACAR 19.19  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.82 1.19 2.26 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 1.98 1.19 2.26 ;
        RECT  0.91 0.82 1.19 1.10 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 32.42  LAYER ME1  ;
        ANTENNADIFFAREA 15.58  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.69  LAYER ME1  ;
        ANTENNAMAXAREACAR 19.19  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.17 1.90 13.45 2.50 ;
        RECT  13.17 0.64 13.45 1.24 ;
        RECT  13.17 0.64 13.33 2.50 ;
        RECT  12.06 1.52 13.33 1.68 ;
        RECT  12.13 1.90 12.41 2.50 ;
        RECT  12.13 0.64 12.41 1.24 ;
        RECT  12.13 0.64 12.34 2.50 ;
        RECT  12.06 1.46 12.34 1.74 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 32.42  LAYER ME1  ;
        ANTENNADIFFAREA 15.61  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.69  LAYER ME1  ;
        ANTENNAMAXAREACAR 19.19  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  15.25 1.90 15.53 2.50 ;
        RECT  15.25 0.64 15.53 1.24 ;
        RECT  15.25 0.64 15.41 2.50 ;
        RECT  14.33 1.52 15.41 1.68 ;
        RECT  14.33 1.46 14.74 1.74 ;
        RECT  14.21 1.90 14.49 2.50 ;
        RECT  14.33 0.64 14.49 2.50 ;
        RECT  14.21 0.64 14.49 1.24 ;
        END
    END QB
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END E
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 16.40 3.48 ;
        RECT  15.83 2.88 16.22 3.48 ;
        RECT  15.77 1.90 16.05 2.50 ;
        RECT  15.83 1.90 15.99 3.48 ;
        RECT  14.73 1.90 15.01 2.50 ;
        RECT  14.79 1.90 14.95 3.48 ;
        RECT  13.69 1.90 13.97 2.50 ;
        RECT  13.75 1.90 13.91 3.48 ;
        RECT  12.65 1.90 12.93 2.50 ;
        RECT  12.71 1.90 12.87 3.48 ;
        RECT  11.61 1.90 11.89 2.50 ;
        RECT  11.67 1.90 11.83 3.48 ;
        RECT  10.37 2.40 10.65 3.48 ;
        RECT  9.57 1.84 9.85 2.12 ;
        RECT  9.63 1.84 9.79 3.48 ;
        RECT  8.57 1.84 8.85 2.12 ;
        RECT  8.63 1.84 8.79 3.48 ;
        RECT  7.57 1.84 7.85 2.12 ;
        RECT  7.67 1.84 7.83 3.48 ;
        RECT  2.71 2.52 2.99 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 16.40 0.28 ;
        RECT  15.83 -0.28 16.22 0.32 ;
        RECT  15.77 0.64 16.05 1.24 ;
        RECT  15.83 -0.28 15.99 1.24 ;
        RECT  14.73 0.64 15.01 1.24 ;
        RECT  14.79 -0.28 14.95 1.24 ;
        RECT  13.69 0.64 13.97 1.24 ;
        RECT  13.75 -0.28 13.91 1.24 ;
        RECT  12.65 0.64 12.93 1.24 ;
        RECT  12.71 -0.28 12.87 1.24 ;
        RECT  11.61 0.64 11.89 1.24 ;
        RECT  11.67 -0.28 11.83 1.24 ;
        RECT  10.61 0.88 10.89 1.16 ;
        RECT  10.67 -0.28 10.83 1.16 ;
        RECT  9.13 -0.28 9.41 0.68 ;
        RECT  2.71 -0.28 2.99 0.64 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.99 0.88 2.27 1.16 ;
        RECT  1.95 1.98 2.23 2.26 ;
        RECT  2.07 0.88 2.23 2.69 ;
        RECT  2.07 2.41 2.37 2.69 ;
        RECT  2.27 0.44 2.55 0.72 ;
        RECT  1.55 0.56 2.55 0.72 ;
        RECT  1.55 0.56 1.71 1.10 ;
        RECT  1.43 0.82 1.71 1.10 ;
        RECT  1.49 0.82 1.65 2.26 ;
        RECT  1.43 1.98 1.71 2.26 ;
        RECT  3.47 0.96 3.86 1.24 ;
        RECT  3.70 1.46 4.02 1.74 ;
        RECT  3.70 0.95 3.86 2.19 ;
        RECT  3.47 1.92 3.75 2.20 ;
        RECT  4.07 0.44 4.35 0.72 ;
        RECT  3.15 0.56 4.35 0.72 ;
        RECT  3.15 0.56 3.31 1.12 ;
        RECT  2.47 0.96 3.31 1.12 ;
        RECT  2.47 0.96 2.75 1.24 ;
        RECT  2.55 0.96 2.71 2.20 ;
        RECT  2.43 1.92 2.71 2.20 ;
        RECT  2.43 2.04 3.31 2.20 ;
        RECT  3.15 2.04 3.31 2.64 ;
        RECT  3.15 2.48 4.25 2.64 ;
        RECT  3.97 2.48 4.25 2.76 ;
        RECT  5.59 0.76 5.91 1.04 ;
        RECT  5.59 0.76 5.75 2.00 ;
        RECT  5.25 1.84 6.29 2.00 ;
        RECT  5.25 1.84 5.53 2.12 ;
        RECT  6.01 1.84 6.29 2.12 ;
        RECT  6.15 0.76 6.43 1.04 ;
        RECT  6.27 0.76 6.43 1.36 ;
        RECT  7.11 1.08 7.39 1.36 ;
        RECT  6.27 1.20 7.39 1.36 ;
        RECT  6.53 1.20 6.69 2.12 ;
        RECT  6.53 1.84 6.81 2.12 ;
        RECT  4.63 0.86 4.91 1.14 ;
        RECT  4.07 0.98 4.91 1.14 ;
        RECT  4.07 0.96 4.35 1.24 ;
        RECT  4.29 0.98 4.45 2.12 ;
        RECT  4.41 1.84 4.57 2.44 ;
        RECT  4.41 2.28 7.51 2.44 ;
        RECT  7.23 2.28 7.51 2.56 ;
        RECT  6.67 0.76 7.95 0.92 ;
        RECT  6.67 0.76 6.95 1.04 ;
        RECT  7.67 0.76 7.95 1.16 ;
        RECT  7.67 0.76 7.83 1.68 ;
        RECT  8.71 1.40 8.99 1.68 ;
        RECT  7.25 1.52 8.99 1.68 ;
        RECT  8.01 1.52 8.17 2.12 ;
        RECT  7.25 1.52 7.41 2.12 ;
        RECT  7.05 1.84 7.41 2.12 ;
        RECT  8.01 1.84 8.37 2.12 ;
        RECT  5.27 0.44 8.87 0.60 ;
        RECT  8.71 0.44 8.87 1.04 ;
        RECT  8.71 0.88 9.37 1.04 ;
        RECT  5.27 0.44 5.43 1.14 ;
        RECT  9.09 0.88 9.37 1.16 ;
        RECT  5.15 0.86 5.31 1.46 ;
        RECT  4.93 1.30 5.31 1.46 ;
        RECT  9.15 0.88 9.31 2.12 ;
        RECT  4.93 1.30 5.09 2.12 ;
        RECT  4.81 1.84 5.09 2.12 ;
        RECT  9.09 1.84 9.37 2.12 ;
        RECT  9.71 0.88 9.99 1.16 ;
        RECT  9.71 1.00 10.27 1.16 ;
        RECT  10.11 1.00 10.27 2.12 ;
        RECT  10.09 1.84 10.37 2.12 ;
        RECT  10.09 1.96 10.97 2.12 ;
        RECT  10.81 1.96 10.97 2.64 ;
        RECT  10.81 2.48 11.44 2.64 ;
        RECT  11.16 2.48 11.44 2.76 ;
        RECT  11.13 0.88 11.41 1.16 ;
        RECT  10.43 1.46 11.55 1.62 ;
        RECT  10.43 1.40 10.71 1.68 ;
        RECT  11.25 1.40 11.55 1.68 ;
        RECT  11.25 0.88 11.41 2.12 ;
        RECT  11.13 1.84 11.41 2.12 ;
    END
END DFFDESSP8V1_0

MACRO DFFDESSP4V1_0
    CLASS CORE ;
    FOREIGN DFFDESSP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 28.14  LAYER ME1  ;
        ANTENNADIFFAREA 12.57  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.11  LAYER ME1  ;
        ANTENNAMAXAREACAR 25.27  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.26 1.46 13.54 1.74 ;
        RECT  13.17 1.90 13.45 2.50 ;
        RECT  13.26 0.64 13.45 2.50 ;
        RECT  13.17 0.64 13.45 1.24 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 28.14  LAYER ME1  ;
        ANTENNADIFFAREA 12.54  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.11  LAYER ME1  ;
        ANTENNAMAXAREACAR 25.27  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.13 1.90 12.41 2.50 ;
        RECT  12.13 0.64 12.41 1.24 ;
        RECT  12.13 0.64 12.34 2.50 ;
        RECT  12.06 1.46 12.34 1.74 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 28.14  LAYER ME1  ;
        ANTENNADIFFAREA 12.45  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.11  LAYER ME1  ;
        ANTENNAMAXAREACAR 25.27  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.82 1.19 2.26 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 1.98 1.19 2.26 ;
        RECT  0.91 0.82 1.19 1.10 ;
        END
    END D
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.53 1.40 9.95 1.68 ;
        END
    END SB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.24 1.40 3.54 1.76 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END E
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 14.40 0.28 ;
        RECT  13.78 -0.28 14.22 0.32 ;
        RECT  13.69 0.64 13.97 1.24 ;
        RECT  13.78 -0.28 13.94 1.24 ;
        RECT  12.65 0.64 12.93 1.24 ;
        RECT  12.71 -0.28 12.87 1.24 ;
        RECT  11.61 0.64 11.89 1.24 ;
        RECT  11.67 -0.28 11.83 1.24 ;
        RECT  10.61 0.88 10.89 1.16 ;
        RECT  10.67 -0.28 10.83 1.16 ;
        RECT  9.13 -0.28 9.41 0.68 ;
        RECT  2.71 -0.28 2.99 0.64 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 14.40 3.48 ;
        RECT  13.78 2.88 14.22 3.48 ;
        RECT  13.69 1.90 13.97 2.50 ;
        RECT  13.78 1.90 13.94 3.48 ;
        RECT  12.65 1.90 12.93 2.50 ;
        RECT  12.71 1.90 12.87 3.48 ;
        RECT  11.61 1.90 11.89 2.50 ;
        RECT  11.67 1.90 11.83 3.48 ;
        RECT  10.37 2.40 10.65 3.48 ;
        RECT  9.57 1.84 9.85 2.12 ;
        RECT  9.63 1.84 9.79 3.48 ;
        RECT  8.57 1.84 8.85 2.12 ;
        RECT  8.63 1.84 8.79 3.48 ;
        RECT  7.57 1.84 7.85 2.12 ;
        RECT  7.67 1.84 7.83 3.48 ;
        RECT  2.71 2.52 2.99 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.99 0.88 2.27 1.16 ;
        RECT  1.95 1.98 2.23 2.26 ;
        RECT  2.07 0.88 2.23 2.69 ;
        RECT  2.07 2.41 2.37 2.69 ;
        RECT  2.27 0.44 2.55 0.72 ;
        RECT  1.55 0.56 2.55 0.72 ;
        RECT  1.55 0.56 1.71 1.10 ;
        RECT  1.43 0.82 1.71 1.10 ;
        RECT  1.49 0.82 1.65 2.26 ;
        RECT  1.43 1.98 1.71 2.26 ;
        RECT  3.47 0.96 3.86 1.24 ;
        RECT  3.70 1.46 4.02 1.74 ;
        RECT  3.70 0.96 3.86 2.20 ;
        RECT  3.47 1.92 3.86 2.20 ;
        RECT  4.07 0.44 4.35 0.72 ;
        RECT  3.15 0.56 4.35 0.72 ;
        RECT  3.15 0.56 3.31 1.12 ;
        RECT  2.47 0.96 3.31 1.12 ;
        RECT  2.47 0.96 2.75 1.24 ;
        RECT  2.55 0.96 2.71 2.20 ;
        RECT  2.43 1.92 2.71 2.20 ;
        RECT  2.43 2.04 3.31 2.20 ;
        RECT  3.15 2.04 3.31 2.64 ;
        RECT  3.15 2.48 4.25 2.64 ;
        RECT  3.97 2.48 4.25 2.76 ;
        RECT  5.59 0.76 5.91 1.04 ;
        RECT  5.59 0.76 5.75 2.00 ;
        RECT  5.25 1.84 6.29 2.00 ;
        RECT  5.25 1.84 5.53 2.12 ;
        RECT  6.01 1.84 6.29 2.12 ;
        RECT  6.15 0.76 6.43 1.04 ;
        RECT  6.27 0.76 6.43 1.36 ;
        RECT  7.11 1.08 7.39 1.36 ;
        RECT  6.27 1.20 7.39 1.36 ;
        RECT  6.53 1.20 6.69 2.12 ;
        RECT  6.53 1.84 6.81 2.12 ;
        RECT  4.63 0.86 4.91 1.14 ;
        RECT  4.07 0.98 4.91 1.14 ;
        RECT  4.07 0.96 4.35 1.24 ;
        RECT  4.29 0.98 4.45 2.12 ;
        RECT  4.41 1.84 4.57 2.44 ;
        RECT  4.41 2.28 7.51 2.44 ;
        RECT  7.23 2.28 7.51 2.56 ;
        RECT  6.67 0.76 7.95 0.92 ;
        RECT  6.67 0.76 6.95 1.04 ;
        RECT  7.67 0.76 7.95 1.16 ;
        RECT  7.67 0.76 7.83 1.68 ;
        RECT  8.71 1.40 8.99 1.68 ;
        RECT  7.25 1.52 8.99 1.68 ;
        RECT  8.01 1.52 8.17 2.12 ;
        RECT  7.25 1.52 7.41 2.12 ;
        RECT  7.05 1.84 7.41 2.12 ;
        RECT  8.01 1.84 8.37 2.12 ;
        RECT  5.27 0.44 8.87 0.60 ;
        RECT  8.71 0.44 8.87 1.04 ;
        RECT  8.71 0.88 9.37 1.04 ;
        RECT  5.27 0.44 5.43 1.14 ;
        RECT  9.09 0.88 9.37 1.16 ;
        RECT  5.15 0.86 5.31 1.46 ;
        RECT  4.93 1.30 5.31 1.46 ;
        RECT  9.15 0.88 9.31 2.12 ;
        RECT  4.93 1.30 5.09 2.12 ;
        RECT  4.81 1.84 5.09 2.12 ;
        RECT  9.09 1.84 9.37 2.12 ;
        RECT  9.71 0.88 9.99 1.16 ;
        RECT  9.71 1.00 10.27 1.16 ;
        RECT  10.11 1.00 10.27 2.12 ;
        RECT  10.09 1.84 10.37 2.12 ;
        RECT  10.09 1.96 10.97 2.12 ;
        RECT  10.81 1.96 10.97 2.64 ;
        RECT  10.81 2.48 11.44 2.64 ;
        RECT  11.16 2.48 11.44 2.76 ;
        RECT  11.13 0.88 11.41 1.16 ;
        RECT  10.43 1.46 11.55 1.62 ;
        RECT  10.43 1.40 10.71 1.68 ;
        RECT  11.25 1.40 11.55 1.68 ;
        RECT  11.25 0.88 11.41 2.12 ;
        RECT  11.13 1.84 11.41 2.12 ;
    END
END DFFDESSP4V1_0

MACRO DFFDESSP2V1_0
    CLASS CORE ;
    FOREIGN DFFDESSP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 13.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.24 1.40 3.54 1.76 ;
        END
    END CK
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.53 1.40 9.95 1.68 ;
        END
    END SB
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 25.95  LAYER ME1  ;
        ANTENNADIFFAREA 11.10  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.83  LAYER ME1  ;
        ANTENNAMAXAREACAR 31.43  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.82 1.19 2.26 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 1.98 1.19 2.26 ;
        RECT  0.91 0.82 1.19 1.10 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 25.95  LAYER ME1  ;
        ANTENNADIFFAREA 10.99  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.83  LAYER ME1  ;
        ANTENNAMAXAREACAR 31.43  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.73 1.46 12.34 1.74 ;
        RECT  11.61 1.90 11.89 2.50 ;
        RECT  11.73 0.64 11.89 2.50 ;
        RECT  11.61 0.64 11.89 1.24 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 25.95  LAYER ME1  ;
        ANTENNADIFFAREA 10.99  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.83  LAYER ME1  ;
        ANTENNAMAXAREACAR 31.43  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.77 1.46 13.12 1.74 ;
        RECT  12.65 1.90 12.93 2.50 ;
        RECT  12.77 0.64 12.93 2.50 ;
        RECT  12.65 0.64 12.93 1.24 ;
        END
    END QB
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END E
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 13.20 3.48 ;
        RECT  12.74 2.88 13.02 3.48 ;
        RECT  12.13 1.90 12.41 2.50 ;
        RECT  12.19 1.90 12.35 3.48 ;
        RECT  10.37 2.40 10.65 3.48 ;
        RECT  9.57 1.84 9.85 2.12 ;
        RECT  9.63 1.84 9.79 3.48 ;
        RECT  8.57 1.84 8.85 2.12 ;
        RECT  8.63 1.84 8.79 3.48 ;
        RECT  7.57 1.84 7.85 2.12 ;
        RECT  7.67 1.84 7.83 3.48 ;
        RECT  2.71 2.52 2.99 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 13.20 0.28 ;
        RECT  12.74 -0.28 13.02 0.32 ;
        RECT  12.13 0.64 12.41 1.24 ;
        RECT  12.19 -0.28 12.35 1.24 ;
        RECT  10.61 0.88 10.89 1.16 ;
        RECT  10.67 -0.28 10.83 1.16 ;
        RECT  9.13 -0.28 9.41 0.68 ;
        RECT  2.71 -0.28 2.99 0.64 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.99 0.88 2.27 1.16 ;
        RECT  1.95 1.98 2.23 2.26 ;
        RECT  2.07 0.88 2.23 2.69 ;
        RECT  2.07 2.41 2.37 2.69 ;
        RECT  2.23 0.44 2.51 0.72 ;
        RECT  1.55 0.56 2.51 0.72 ;
        RECT  1.55 0.56 1.71 1.10 ;
        RECT  1.43 0.82 1.71 1.10 ;
        RECT  1.49 0.82 1.65 2.26 ;
        RECT  1.43 1.98 1.71 2.26 ;
        RECT  3.47 0.96 3.86 1.24 ;
        RECT  3.70 1.46 4.02 1.74 ;
        RECT  3.70 0.96 3.86 2.20 ;
        RECT  3.47 1.92 3.86 2.20 ;
        RECT  4.07 0.44 4.35 0.72 ;
        RECT  3.15 0.56 4.35 0.72 ;
        RECT  3.15 0.56 3.31 1.12 ;
        RECT  2.47 0.96 3.31 1.12 ;
        RECT  2.47 0.96 2.75 1.24 ;
        RECT  2.55 0.96 2.71 2.20 ;
        RECT  2.43 1.92 2.71 2.20 ;
        RECT  2.43 2.04 3.31 2.20 ;
        RECT  3.15 2.04 3.31 2.64 ;
        RECT  3.15 2.48 4.25 2.64 ;
        RECT  3.97 2.48 4.25 2.76 ;
        RECT  5.59 0.76 5.91 1.04 ;
        RECT  5.59 0.76 5.75 2.00 ;
        RECT  5.25 1.84 6.29 2.00 ;
        RECT  5.25 1.84 5.53 2.12 ;
        RECT  6.01 1.84 6.29 2.12 ;
        RECT  6.15 0.76 6.43 1.04 ;
        RECT  6.27 0.76 6.43 1.36 ;
        RECT  7.11 1.08 7.39 1.36 ;
        RECT  6.27 1.20 7.39 1.36 ;
        RECT  6.53 1.20 6.69 2.12 ;
        RECT  6.53 1.84 6.81 2.12 ;
        RECT  4.63 0.86 4.91 1.14 ;
        RECT  4.07 0.98 4.91 1.14 ;
        RECT  4.07 0.96 4.35 1.24 ;
        RECT  4.29 0.98 4.45 2.12 ;
        RECT  4.41 1.84 4.57 2.44 ;
        RECT  4.41 2.28 7.51 2.44 ;
        RECT  7.23 2.28 7.51 2.56 ;
        RECT  6.67 0.76 7.95 0.92 ;
        RECT  6.67 0.76 6.95 1.04 ;
        RECT  7.67 0.76 7.95 1.16 ;
        RECT  7.67 0.76 7.83 1.68 ;
        RECT  8.71 1.40 8.99 1.68 ;
        RECT  7.25 1.52 8.99 1.68 ;
        RECT  8.01 1.52 8.17 2.12 ;
        RECT  7.25 1.52 7.41 2.12 ;
        RECT  7.05 1.84 7.41 2.12 ;
        RECT  8.01 1.84 8.37 2.12 ;
        RECT  5.27 0.44 8.87 0.60 ;
        RECT  8.71 0.44 8.87 1.04 ;
        RECT  8.71 0.88 9.37 1.04 ;
        RECT  5.27 0.44 5.43 1.14 ;
        RECT  9.09 0.88 9.37 1.16 ;
        RECT  5.15 0.86 5.31 1.46 ;
        RECT  4.93 1.30 5.31 1.46 ;
        RECT  9.15 0.88 9.31 2.12 ;
        RECT  4.93 1.30 5.09 2.12 ;
        RECT  4.81 1.84 5.09 2.12 ;
        RECT  9.09 1.84 9.37 2.12 ;
        RECT  9.71 0.88 9.99 1.16 ;
        RECT  9.71 1.00 10.27 1.16 ;
        RECT  10.11 1.00 10.27 2.12 ;
        RECT  10.09 1.84 10.37 2.12 ;
        RECT  10.09 1.96 10.97 2.12 ;
        RECT  10.81 1.96 10.97 2.64 ;
        RECT  10.81 2.48 11.44 2.64 ;
        RECT  11.16 2.48 11.44 2.76 ;
        RECT  11.13 0.88 11.41 1.16 ;
        RECT  10.43 1.46 11.55 1.62 ;
        RECT  10.43 1.40 10.71 1.68 ;
        RECT  11.25 1.40 11.55 1.68 ;
        RECT  11.25 0.88 11.41 2.12 ;
        RECT  11.13 1.84 11.41 2.12 ;
    END
END DFFDESSP2V1_0

MACRO DFFDESSP1V1_0
    CLASS CORE ;
    FOREIGN DFFDESSP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 13.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 25.50  LAYER ME1  ;
        ANTENNADIFFAREA 10.41  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER ME1  ;
        ANTENNAMAXAREACAR 37.95  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.82 1.19 2.26 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 1.98 1.19 2.26 ;
        RECT  0.91 0.82 1.19 1.10 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 25.50  LAYER ME1  ;
        ANTENNADIFFAREA 10.30  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER ME1  ;
        ANTENNAMAXAREACAR 37.95  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.73 1.46 12.34 1.74 ;
        RECT  11.61 1.90 11.89 2.18 ;
        RECT  11.73 0.96 11.89 2.18 ;
        RECT  11.61 0.96 11.89 1.24 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.53 1.40 9.95 1.68 ;
        END
    END SB
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 25.19  LAYER ME1  ;
        ANTENNADIFFAREA 10.30  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER ME1  ;
        ANTENNAMAXAREACAR 37.48  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.77 1.46 13.12 1.74 ;
        RECT  12.65 1.90 12.93 2.18 ;
        RECT  12.77 0.96 12.93 2.18 ;
        RECT  12.65 0.96 12.93 1.24 ;
        END
    END QB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.24 1.40 3.54 1.76 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END E
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 13.20 3.48 ;
        RECT  12.74 2.88 13.02 3.48 ;
        RECT  12.13 1.90 12.41 2.18 ;
        RECT  12.19 1.90 12.35 3.48 ;
        RECT  10.37 2.40 10.65 3.48 ;
        RECT  9.57 1.84 9.85 2.12 ;
        RECT  9.63 1.84 9.79 3.48 ;
        RECT  8.57 1.84 8.85 2.12 ;
        RECT  8.63 1.84 8.79 3.48 ;
        RECT  7.57 1.84 7.85 2.12 ;
        RECT  7.67 1.84 7.83 3.48 ;
        RECT  2.71 2.52 2.99 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 13.20 0.28 ;
        RECT  12.74 -0.28 13.02 0.32 ;
        RECT  12.13 0.96 12.41 1.24 ;
        RECT  12.19 -0.28 12.35 1.24 ;
        RECT  10.61 0.88 10.89 1.16 ;
        RECT  10.67 -0.28 10.83 1.16 ;
        RECT  9.13 -0.28 9.41 0.68 ;
        RECT  2.71 -0.28 2.99 0.64 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.99 0.88 2.27 1.16 ;
        RECT  1.95 1.98 2.23 2.26 ;
        RECT  2.07 0.88 2.23 2.70 ;
        RECT  2.07 2.42 2.37 2.70 ;
        RECT  1.55 0.50 2.37 0.66 ;
        RECT  2.09 0.44 2.37 0.72 ;
        RECT  1.55 0.50 1.71 1.10 ;
        RECT  1.43 0.82 1.71 1.10 ;
        RECT  1.49 0.82 1.65 2.26 ;
        RECT  1.43 1.98 1.71 2.26 ;
        RECT  3.47 0.96 3.86 1.24 ;
        RECT  3.70 1.46 4.02 1.74 ;
        RECT  3.70 0.96 3.86 2.20 ;
        RECT  3.47 1.92 3.86 2.20 ;
        RECT  4.07 0.44 4.35 0.72 ;
        RECT  3.15 0.56 4.35 0.72 ;
        RECT  3.15 0.56 3.31 1.12 ;
        RECT  2.47 0.96 3.31 1.12 ;
        RECT  2.47 0.96 2.75 1.24 ;
        RECT  2.55 0.96 2.71 2.20 ;
        RECT  2.43 1.92 2.71 2.20 ;
        RECT  2.43 2.04 3.31 2.20 ;
        RECT  3.15 2.04 3.31 2.64 ;
        RECT  3.15 2.48 4.25 2.64 ;
        RECT  3.97 2.48 4.25 2.76 ;
        RECT  5.59 0.76 5.91 1.04 ;
        RECT  5.59 0.76 5.75 2.00 ;
        RECT  5.25 1.84 6.29 2.00 ;
        RECT  5.25 1.84 5.53 2.12 ;
        RECT  6.01 1.84 6.29 2.12 ;
        RECT  6.15 0.76 6.43 1.04 ;
        RECT  6.27 0.76 6.43 1.36 ;
        RECT  7.11 1.08 7.39 1.36 ;
        RECT  6.27 1.20 7.39 1.36 ;
        RECT  6.53 1.20 6.69 2.12 ;
        RECT  6.53 1.84 6.81 2.12 ;
        RECT  4.63 0.86 4.91 1.14 ;
        RECT  4.07 0.98 4.91 1.14 ;
        RECT  4.07 0.96 4.35 1.24 ;
        RECT  4.29 0.98 4.45 2.12 ;
        RECT  4.41 1.84 4.57 2.44 ;
        RECT  4.41 2.28 7.51 2.44 ;
        RECT  7.23 2.28 7.51 2.56 ;
        RECT  6.67 0.76 7.95 0.92 ;
        RECT  6.67 0.76 6.95 1.04 ;
        RECT  7.67 0.76 7.95 1.16 ;
        RECT  7.67 0.76 7.83 1.68 ;
        RECT  8.71 1.40 8.99 1.68 ;
        RECT  7.25 1.52 8.99 1.68 ;
        RECT  8.01 1.52 8.17 2.12 ;
        RECT  7.25 1.52 7.41 2.12 ;
        RECT  7.05 1.84 7.41 2.12 ;
        RECT  8.01 1.84 8.37 2.12 ;
        RECT  5.27 0.44 8.87 0.60 ;
        RECT  8.71 0.44 8.87 1.04 ;
        RECT  8.71 0.88 9.37 1.04 ;
        RECT  5.27 0.44 5.43 1.14 ;
        RECT  9.09 0.88 9.37 1.16 ;
        RECT  5.15 0.86 5.31 1.46 ;
        RECT  4.93 1.30 5.31 1.46 ;
        RECT  9.15 0.88 9.31 2.12 ;
        RECT  4.93 1.30 5.09 2.12 ;
        RECT  4.81 1.84 5.09 2.12 ;
        RECT  9.09 1.84 9.37 2.12 ;
        RECT  9.71 0.88 9.99 1.16 ;
        RECT  9.71 1.00 10.27 1.16 ;
        RECT  10.11 1.00 10.27 2.12 ;
        RECT  10.09 1.84 10.37 2.12 ;
        RECT  10.09 1.96 10.97 2.12 ;
        RECT  10.81 1.96 10.97 2.64 ;
        RECT  10.81 2.48 11.44 2.64 ;
        RECT  11.16 2.48 11.44 2.76 ;
        RECT  11.13 0.88 11.41 1.16 ;
        RECT  10.43 1.46 11.55 1.62 ;
        RECT  10.43 1.40 10.71 1.68 ;
        RECT  11.25 1.40 11.55 1.68 ;
        RECT  11.25 0.88 11.41 2.12 ;
        RECT  11.13 1.84 11.41 2.12 ;
    END
END DFFDESSP1V1_0

MACRO DFFDESP8V1_0
    CLASS CORE ;
    FOREIGN DFFDESP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 25.98  LAYER ME1  ;
        ANTENNADIFFAREA 12.98  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.69  LAYER ME1  ;
        ANTENNAMAXAREACAR 15.38  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.97 1.90 13.25 2.18 ;
        RECT  12.97 0.96 13.25 1.24 ;
        RECT  12.97 0.96 13.13 2.18 ;
        RECT  12.05 1.52 13.13 1.68 ;
        RECT  12.05 1.46 12.34 1.74 ;
        RECT  11.93 1.90 12.21 2.18 ;
        RECT  12.05 0.96 12.21 2.18 ;
        RECT  11.93 0.96 12.21 1.24 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 25.98  LAYER ME1  ;
        ANTENNADIFFAREA 12.98  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.69  LAYER ME1  ;
        ANTENNAMAXAREACAR 15.38  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.89 1.90 11.17 2.18 ;
        RECT  10.89 0.96 11.17 1.24 ;
        RECT  10.89 0.96 11.05 2.18 ;
        RECT  9.97 1.52 11.05 1.68 ;
        RECT  9.97 1.46 10.34 1.74 ;
        RECT  9.85 1.90 10.13 2.18 ;
        RECT  9.97 0.96 10.13 2.18 ;
        RECT  9.85 0.96 10.13 1.24 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 25.98  LAYER ME1  ;
        ANTENNADIFFAREA 12.89  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.69  LAYER ME1  ;
        ANTENNAMAXAREACAR 15.38  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.81 1.19 2.25 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  0.91 0.81 1.19 1.09 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.87 1.46 3.37 1.74 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END E
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 14.00 0.28 ;
        RECT  13.54 -0.28 13.82 0.32 ;
        RECT  13.49 0.64 13.77 0.92 ;
        RECT  13.55 -0.28 13.71 0.92 ;
        RECT  12.45 0.64 12.73 0.92 ;
        RECT  12.51 -0.28 12.67 0.92 ;
        RECT  11.41 0.64 11.69 0.92 ;
        RECT  11.47 -0.28 11.63 0.92 ;
        RECT  10.37 0.64 10.65 0.92 ;
        RECT  10.43 -0.28 10.59 0.92 ;
        RECT  9.33 0.64 9.61 0.92 ;
        RECT  9.39 -0.28 9.55 0.92 ;
        RECT  8.33 0.96 8.61 1.24 ;
        RECT  8.43 -0.28 8.59 1.24 ;
        RECT  5.59 0.72 5.87 1.00 ;
        RECT  5.65 -0.28 5.81 1.00 ;
        RECT  2.95 0.88 3.23 1.16 ;
        RECT  3.05 -0.28 3.21 1.16 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 14.00 3.48 ;
        RECT  13.54 2.88 13.82 3.48 ;
        RECT  13.49 2.22 13.77 2.50 ;
        RECT  13.55 2.22 13.71 3.48 ;
        RECT  12.45 2.22 12.73 2.50 ;
        RECT  12.51 2.22 12.67 3.48 ;
        RECT  11.41 2.22 11.69 2.50 ;
        RECT  11.47 2.22 11.63 3.48 ;
        RECT  10.37 2.22 10.65 2.50 ;
        RECT  10.43 2.22 10.59 3.48 ;
        RECT  9.33 2.22 9.61 2.50 ;
        RECT  9.39 2.22 9.55 3.48 ;
        RECT  8.33 1.84 8.61 2.12 ;
        RECT  8.39 1.84 8.55 3.48 ;
        RECT  5.77 1.92 6.05 2.20 ;
        RECT  5.83 1.92 5.99 3.48 ;
        RECT  2.74 2.52 3.02 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.95 0.81 2.23 1.09 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.81 2.23 2.63 ;
        RECT  2.07 2.35 2.37 2.63 ;
        RECT  1.55 0.49 2.89 0.65 ;
        RECT  2.61 0.44 2.89 0.72 ;
        RECT  1.55 0.49 1.71 1.09 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  3.47 0.88 3.77 1.16 ;
        RECT  3.61 1.26 3.89 1.54 ;
        RECT  3.61 0.88 3.77 2.14 ;
        RECT  3.49 1.86 3.77 2.14 ;
        RECT  3.97 0.72 4.25 1.00 ;
        RECT  2.43 0.88 2.71 1.16 ;
        RECT  4.05 0.72 4.21 2.20 ;
        RECT  2.55 0.88 2.71 2.14 ;
        RECT  2.43 1.86 2.71 2.14 ;
        RECT  2.43 1.98 3.33 2.14 ;
        RECT  3.97 1.92 4.25 2.20 ;
        RECT  3.17 1.98 3.33 2.46 ;
        RECT  3.97 1.92 4.13 2.46 ;
        RECT  3.17 2.30 4.13 2.46 ;
        RECT  5.05 0.72 5.35 1.00 ;
        RECT  5.05 0.72 5.21 2.20 ;
        RECT  5.01 1.92 5.29 2.20 ;
        RECT  4.49 0.72 4.77 1.00 ;
        RECT  5.85 1.48 6.13 1.76 ;
        RECT  5.45 1.60 6.13 1.76 ;
        RECT  4.55 0.72 4.71 2.20 ;
        RECT  4.49 1.92 4.77 2.20 ;
        RECT  4.61 1.92 4.77 2.52 ;
        RECT  5.45 1.60 5.61 2.52 ;
        RECT  4.61 2.36 5.61 2.52 ;
        RECT  6.11 0.72 6.45 1.00 ;
        RECT  5.37 1.16 6.45 1.32 ;
        RECT  5.37 1.16 5.65 1.44 ;
        RECT  6.29 0.72 6.45 2.20 ;
        RECT  6.29 1.92 6.57 2.20 ;
        RECT  7.19 0.76 7.61 1.04 ;
        RECT  7.33 1.92 7.61 2.20 ;
        RECT  7.45 0.76 7.61 2.76 ;
        RECT  7.45 2.48 7.73 2.76 ;
        RECT  6.79 0.44 8.27 0.60 ;
        RECT  7.99 0.44 8.27 0.80 ;
        RECT  6.67 0.76 6.95 1.04 ;
        RECT  6.79 0.44 6.95 2.20 ;
        RECT  6.79 1.92 7.09 2.20 ;
        RECT  7.81 0.96 8.09 1.24 ;
        RECT  7.81 1.46 8.75 1.62 ;
        RECT  8.47 1.40 8.75 1.68 ;
        RECT  7.81 0.96 7.97 2.12 ;
        RECT  7.81 1.84 8.09 2.12 ;
        RECT  8.85 0.96 9.13 1.24 ;
        RECT  8.85 1.84 9.13 2.12 ;
        RECT  8.97 0.96 9.13 2.76 ;
        RECT  8.88 2.48 9.16 2.76 ;
    END
END DFFDESP8V1_0

MACRO DFFDESP4V1_0
    CLASS CORE ;
    FOREIGN DFFDESP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 22.50  LAYER ME1  ;
        ANTENNADIFFAREA 10.22  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.11  LAYER ME1  ;
        ANTENNAMAXAREACAR 20.21  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.89 1.90 11.17 2.18 ;
        RECT  10.89 0.96 11.17 1.24 ;
        RECT  10.89 0.96 11.14 2.18 ;
        RECT  10.86 1.46 11.14 1.74 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 22.50  LAYER ME1  ;
        ANTENNADIFFAREA 10.22  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.11  LAYER ME1  ;
        ANTENNAMAXAREACAR 20.21  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.97 1.46 10.34 1.74 ;
        RECT  9.85 1.90 10.13 2.18 ;
        RECT  9.97 0.96 10.13 2.18 ;
        RECT  9.85 0.96 10.13 1.24 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.87 1.46 3.37 1.74 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 22.50  LAYER ME1  ;
        ANTENNADIFFAREA 10.33  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.11  LAYER ME1  ;
        ANTENNAMAXAREACAR 20.21  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.81 1.19 2.25 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  0.91 0.81 1.19 1.09 ;
        END
    END D
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 12.00 0.28 ;
        RECT  11.47 -0.28 11.82 0.32 ;
        RECT  11.41 0.64 11.69 0.92 ;
        RECT  11.47 -0.28 11.63 0.92 ;
        RECT  10.37 0.64 10.65 0.92 ;
        RECT  10.43 -0.28 10.59 0.92 ;
        RECT  9.33 0.64 9.61 0.92 ;
        RECT  9.39 -0.28 9.55 0.92 ;
        RECT  8.33 0.96 8.61 1.24 ;
        RECT  8.43 -0.28 8.59 1.24 ;
        RECT  5.59 0.72 5.87 1.00 ;
        RECT  5.65 -0.28 5.81 1.00 ;
        RECT  2.95 0.88 3.23 1.16 ;
        RECT  3.05 -0.28 3.21 1.16 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 12.00 3.48 ;
        RECT  11.47 2.88 11.82 3.48 ;
        RECT  11.41 2.22 11.69 2.50 ;
        RECT  11.47 2.22 11.63 3.48 ;
        RECT  10.37 2.22 10.65 2.50 ;
        RECT  10.43 2.22 10.59 3.48 ;
        RECT  9.33 2.22 9.61 2.50 ;
        RECT  9.39 2.22 9.55 3.48 ;
        RECT  8.33 1.84 8.61 2.12 ;
        RECT  8.39 1.84 8.55 3.48 ;
        RECT  5.77 1.92 6.05 2.20 ;
        RECT  5.83 1.92 5.99 3.48 ;
        RECT  2.74 2.52 3.02 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.95 0.81 2.23 1.09 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.81 2.23 2.63 ;
        RECT  2.07 2.35 2.37 2.63 ;
        RECT  1.55 0.49 2.89 0.65 ;
        RECT  2.61 0.44 2.89 0.72 ;
        RECT  1.55 0.49 1.71 1.09 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  3.47 0.88 3.77 1.16 ;
        RECT  3.61 1.26 3.89 1.54 ;
        RECT  3.61 0.88 3.77 2.14 ;
        RECT  3.49 1.86 3.77 2.14 ;
        RECT  3.97 0.72 4.25 1.00 ;
        RECT  2.43 0.88 2.71 1.16 ;
        RECT  4.05 0.72 4.21 2.20 ;
        RECT  2.55 0.88 2.71 2.14 ;
        RECT  2.43 1.86 2.71 2.14 ;
        RECT  2.43 1.98 3.33 2.14 ;
        RECT  3.97 1.92 4.25 2.20 ;
        RECT  3.17 1.98 3.33 2.46 ;
        RECT  3.97 1.92 4.13 2.46 ;
        RECT  3.17 2.30 4.13 2.46 ;
        RECT  5.05 0.72 5.35 1.00 ;
        RECT  5.05 0.72 5.21 2.20 ;
        RECT  5.01 1.92 5.29 2.20 ;
        RECT  4.49 0.72 4.77 1.00 ;
        RECT  5.85 1.48 6.13 1.76 ;
        RECT  5.45 1.60 6.13 1.76 ;
        RECT  4.55 0.72 4.71 2.20 ;
        RECT  4.49 1.92 4.77 2.20 ;
        RECT  4.61 1.92 4.77 2.52 ;
        RECT  5.45 1.60 5.61 2.52 ;
        RECT  4.61 2.36 5.61 2.52 ;
        RECT  6.11 0.72 6.45 1.00 ;
        RECT  5.37 1.16 6.45 1.32 ;
        RECT  5.37 1.16 5.65 1.44 ;
        RECT  6.29 0.72 6.45 2.20 ;
        RECT  6.29 1.92 6.57 2.20 ;
        RECT  7.19 0.76 7.61 1.04 ;
        RECT  7.33 1.92 7.61 2.20 ;
        RECT  7.45 0.76 7.61 2.76 ;
        RECT  7.45 2.48 7.73 2.76 ;
        RECT  6.79 0.44 8.27 0.60 ;
        RECT  7.99 0.44 8.27 0.80 ;
        RECT  6.67 0.76 6.95 1.04 ;
        RECT  6.79 0.44 6.95 2.20 ;
        RECT  6.79 1.92 7.09 2.20 ;
        RECT  7.81 0.96 8.09 1.24 ;
        RECT  7.81 1.46 8.75 1.62 ;
        RECT  8.47 1.40 8.75 1.68 ;
        RECT  7.81 0.96 7.97 2.12 ;
        RECT  7.81 1.84 8.09 2.12 ;
        RECT  8.85 0.96 9.13 1.24 ;
        RECT  8.85 1.84 9.13 2.12 ;
        RECT  8.97 0.96 9.13 2.76 ;
        RECT  8.88 2.48 9.16 2.76 ;
    END
END DFFDESP4V1_0

MACRO DFFDESP2V1_0
    CLASS CORE ;
    FOREIGN DFFDESP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 20.61  LAYER ME1  ;
        ANTENNADIFFAREA 8.99  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.83  LAYER ME1  ;
        ANTENNAMAXAREACAR 24.96  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.81 1.19 2.25 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  0.91 0.81 1.19 1.09 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.87 1.46 3.37 1.74 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 20.31  LAYER ME1  ;
        ANTENNADIFFAREA 8.99  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.83  LAYER ME1  ;
        ANTENNAMAXAREACAR 24.60  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.46 1.46 10.72 1.74 ;
        RECT  10.37 1.90 10.65 2.18 ;
        RECT  10.46 0.96 10.65 2.18 ;
        RECT  10.37 0.96 10.65 1.24 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 20.61  LAYER ME1  ;
        ANTENNADIFFAREA 8.99  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.83  LAYER ME1  ;
        ANTENNAMAXAREACAR 24.96  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.45 1.46 9.94 1.74 ;
        RECT  9.33 1.90 9.61 2.18 ;
        RECT  9.45 0.96 9.61 2.18 ;
        RECT  9.33 0.96 9.61 1.24 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END E
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 10.80 3.48 ;
        RECT  10.34 2.88 10.62 3.48 ;
        RECT  9.85 2.22 10.13 2.50 ;
        RECT  9.91 2.22 10.07 3.48 ;
        RECT  8.33 1.84 8.61 2.12 ;
        RECT  8.39 1.84 8.55 3.48 ;
        RECT  5.77 1.92 6.05 2.20 ;
        RECT  5.83 1.92 5.99 3.48 ;
        RECT  2.74 2.52 3.02 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 10.80 0.28 ;
        RECT  10.34 -0.28 10.62 0.32 ;
        RECT  9.85 0.64 10.13 0.92 ;
        RECT  9.91 -0.28 10.07 0.92 ;
        RECT  8.33 0.96 8.61 1.24 ;
        RECT  8.43 -0.28 8.59 1.24 ;
        RECT  5.59 0.72 5.87 1.00 ;
        RECT  5.65 -0.28 5.81 1.00 ;
        RECT  2.95 0.88 3.23 1.16 ;
        RECT  3.05 -0.28 3.21 1.16 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.95 0.81 2.23 1.09 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.81 2.23 2.63 ;
        RECT  2.07 2.35 2.37 2.63 ;
        RECT  1.55 0.49 2.89 0.65 ;
        RECT  2.61 0.44 2.89 0.72 ;
        RECT  1.55 0.49 1.71 1.09 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  3.47 0.88 3.77 1.16 ;
        RECT  3.61 1.26 3.89 1.54 ;
        RECT  3.61 0.88 3.77 2.14 ;
        RECT  3.49 1.86 3.77 2.14 ;
        RECT  3.97 0.72 4.25 1.00 ;
        RECT  2.43 0.88 2.71 1.16 ;
        RECT  4.05 0.72 4.21 2.20 ;
        RECT  2.55 0.88 2.71 2.14 ;
        RECT  2.43 1.86 2.71 2.14 ;
        RECT  2.43 1.98 3.33 2.14 ;
        RECT  3.97 1.92 4.25 2.20 ;
        RECT  3.17 1.98 3.33 2.46 ;
        RECT  3.97 1.92 4.13 2.46 ;
        RECT  3.17 2.30 4.13 2.46 ;
        RECT  5.05 0.72 5.35 1.00 ;
        RECT  5.05 0.72 5.21 2.20 ;
        RECT  5.01 1.92 5.29 2.20 ;
        RECT  4.49 0.72 4.77 1.00 ;
        RECT  5.85 1.48 6.13 1.76 ;
        RECT  5.45 1.60 6.13 1.76 ;
        RECT  4.55 0.72 4.71 2.20 ;
        RECT  4.49 1.92 4.77 2.20 ;
        RECT  4.61 1.92 4.77 2.52 ;
        RECT  5.45 1.60 5.61 2.52 ;
        RECT  4.61 2.36 5.61 2.52 ;
        RECT  6.11 0.72 6.45 1.00 ;
        RECT  5.37 1.16 6.45 1.32 ;
        RECT  5.37 1.16 5.65 1.44 ;
        RECT  6.29 0.72 6.45 2.20 ;
        RECT  6.29 1.92 6.57 2.20 ;
        RECT  7.19 0.76 7.61 1.04 ;
        RECT  7.33 1.92 7.61 2.20 ;
        RECT  7.45 0.76 7.61 2.76 ;
        RECT  7.45 2.48 7.73 2.76 ;
        RECT  6.79 0.44 8.27 0.60 ;
        RECT  7.99 0.44 8.27 0.80 ;
        RECT  6.67 0.76 6.95 1.04 ;
        RECT  6.79 0.44 6.95 2.20 ;
        RECT  6.79 1.92 7.09 2.20 ;
        RECT  7.81 0.96 8.09 1.24 ;
        RECT  7.81 1.46 8.75 1.62 ;
        RECT  8.47 1.40 8.75 1.68 ;
        RECT  7.81 0.96 7.97 2.12 ;
        RECT  7.81 1.84 8.09 2.12 ;
        RECT  8.85 0.96 9.13 1.24 ;
        RECT  8.85 1.84 9.13 2.12 ;
        RECT  8.97 0.96 9.13 2.76 ;
        RECT  8.88 2.48 9.16 2.76 ;
    END
END DFFDESP2V1_0

MACRO DFFDESP1V1_0
    CLASS CORE ;
    FOREIGN DFFDESP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 20.39  LAYER ME1  ;
        ANTENNADIFFAREA 8.18  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER ME1  ;
        ANTENNAMAXAREACAR 30.35  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.33 1.90 9.61 2.18 ;
        RECT  9.33 0.96 9.61 1.24 ;
        RECT  9.26 1.46 9.54 1.74 ;
        RECT  9.33 0.96 9.49 2.18 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 20.69  LAYER ME1  ;
        ANTENNADIFFAREA 8.18  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER ME1  ;
        ANTENNAMAXAREACAR 30.79  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.37 1.90 10.65 2.18 ;
        RECT  10.37 0.96 10.65 1.24 ;
        RECT  10.37 0.96 10.53 2.18 ;
        RECT  10.06 1.46 10.53 1.74 ;
        END
    END QB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.87 1.46 3.37 1.74 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 20.69  LAYER ME1  ;
        ANTENNADIFFAREA 8.29  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER ME1  ;
        ANTENNAMAXAREACAR 30.79  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.81 1.19 2.25 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  0.91 0.81 1.19 1.09 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END E
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 10.80 0.28 ;
        RECT  10.34 -0.28 10.62 0.32 ;
        RECT  9.85 0.96 10.13 1.24 ;
        RECT  9.91 -0.28 10.07 1.24 ;
        RECT  8.33 0.96 8.61 1.24 ;
        RECT  8.43 -0.28 8.59 1.24 ;
        RECT  5.59 0.72 5.87 1.00 ;
        RECT  5.65 -0.28 5.81 1.00 ;
        RECT  2.95 0.88 3.23 1.16 ;
        RECT  3.05 -0.28 3.21 1.16 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 10.80 3.48 ;
        RECT  10.34 2.88 10.62 3.48 ;
        RECT  9.85 1.90 10.13 2.18 ;
        RECT  9.91 1.90 10.07 3.48 ;
        RECT  8.33 1.84 8.61 2.12 ;
        RECT  8.39 1.84 8.55 3.48 ;
        RECT  5.77 1.92 6.05 2.20 ;
        RECT  5.83 1.92 5.99 3.48 ;
        RECT  2.74 2.52 3.02 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.95 0.81 2.23 1.09 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.81 2.23 2.63 ;
        RECT  2.07 2.35 2.37 2.63 ;
        RECT  1.55 0.49 2.89 0.65 ;
        RECT  2.61 0.44 2.89 0.72 ;
        RECT  1.55 0.49 1.71 1.09 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  3.47 0.88 3.77 1.16 ;
        RECT  3.61 1.26 3.89 1.54 ;
        RECT  3.61 0.88 3.77 2.14 ;
        RECT  3.49 1.86 3.77 2.14 ;
        RECT  3.97 0.72 4.25 1.00 ;
        RECT  2.43 0.88 2.71 1.16 ;
        RECT  4.05 0.72 4.21 2.20 ;
        RECT  2.55 0.88 2.71 2.14 ;
        RECT  2.43 1.86 2.71 2.14 ;
        RECT  2.43 1.98 3.33 2.14 ;
        RECT  3.97 1.92 4.25 2.20 ;
        RECT  3.17 1.98 3.33 2.46 ;
        RECT  3.97 1.92 4.13 2.46 ;
        RECT  3.17 2.30 4.13 2.46 ;
        RECT  5.05 0.72 5.35 1.00 ;
        RECT  5.05 0.72 5.21 2.20 ;
        RECT  5.01 1.92 5.29 2.20 ;
        RECT  4.49 0.72 4.77 1.00 ;
        RECT  5.85 1.48 6.13 1.76 ;
        RECT  5.45 1.60 6.13 1.76 ;
        RECT  4.55 0.72 4.71 2.20 ;
        RECT  4.49 1.92 4.77 2.20 ;
        RECT  4.61 1.92 4.77 2.52 ;
        RECT  5.45 1.60 5.61 2.52 ;
        RECT  4.61 2.36 5.61 2.52 ;
        RECT  6.11 0.72 6.45 1.00 ;
        RECT  5.37 1.16 6.45 1.32 ;
        RECT  5.37 1.16 5.65 1.44 ;
        RECT  6.29 0.72 6.45 2.20 ;
        RECT  6.29 1.92 6.57 2.20 ;
        RECT  7.19 0.76 7.61 1.04 ;
        RECT  7.33 1.92 7.61 2.20 ;
        RECT  7.45 0.76 7.61 2.70 ;
        RECT  7.45 2.42 7.75 2.70 ;
        RECT  6.79 0.44 8.27 0.60 ;
        RECT  7.99 0.44 8.27 0.80 ;
        RECT  6.67 0.76 6.95 1.04 ;
        RECT  6.79 0.44 6.95 2.20 ;
        RECT  6.79 1.92 7.09 2.20 ;
        RECT  7.81 0.96 8.09 1.24 ;
        RECT  7.81 1.46 8.75 1.62 ;
        RECT  8.47 1.40 8.75 1.68 ;
        RECT  7.81 0.96 7.97 2.12 ;
        RECT  7.81 1.84 8.09 2.12 ;
        RECT  8.85 0.96 9.13 1.24 ;
        RECT  8.85 1.84 9.13 2.12 ;
        RECT  8.94 0.96 9.10 2.70 ;
        RECT  8.94 2.42 9.23 2.70 ;
    END
END DFFDESP1V1_0

MACRO DFFDERZSP8V1_0
    CLASS CORE ;
    FOREIGN DFFDERZSP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 36.18  LAYER ME1  ;
        ANTENNADIFFAREA 17.42  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.76  LAYER ME1  ;
        ANTENNAMAXAREACAR 20.59  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  17.26 1.90 17.54 2.50 ;
        RECT  17.26 0.64 17.54 1.24 ;
        RECT  17.26 0.64 17.42 2.50 ;
        RECT  16.34 1.52 17.42 1.68 ;
        RECT  16.34 1.46 16.74 1.74 ;
        RECT  16.22 1.90 16.50 2.50 ;
        RECT  16.34 0.64 16.50 2.50 ;
        RECT  16.22 0.64 16.50 1.24 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 36.18  LAYER ME1  ;
        ANTENNADIFFAREA 17.17  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.76  LAYER ME1  ;
        ANTENNAMAXAREACAR 20.59  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  15.18 1.90 15.46 2.50 ;
        RECT  15.18 0.64 15.46 1.24 ;
        RECT  15.18 0.64 15.34 2.50 ;
        RECT  14.06 1.52 15.34 1.68 ;
        RECT  14.14 1.90 14.42 2.50 ;
        RECT  14.14 0.64 14.42 1.24 ;
        RECT  14.14 0.64 14.34 2.50 ;
        RECT  14.06 1.46 14.34 1.74 ;
        END
    END Q
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.57 1.40 11.95 1.68 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.63 1.40 5.94 1.76 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 36.18  LAYER ME1  ;
        ANTENNADIFFAREA 16.70  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.76  LAYER ME1  ;
        ANTENNAMAXAREACAR 20.59  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.42 1.46 4.74 1.74 ;
        RECT  4.34 0.88 4.62 1.16 ;
        RECT  4.30 1.98 4.58 2.26 ;
        RECT  4.42 0.88 4.58 2.26 ;
        END
    END TD
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 35.86  LAYER ME1  ;
        ANTENNADIFFAREA 16.70  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.76  LAYER ME1  ;
        ANTENNAMAXAREACAR 20.41  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.21 1.88 1.51 2.16 ;
        RECT  1.21 0.66 1.51 0.96 ;
        RECT  1.21 0.66 1.37 2.16 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.99 1.46 2.34 1.76 ;
        END
    END E
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.45 1.06 2.78 1.34 ;
        RECT  2.26 1.06 2.78 1.30 ;
        END
    END SEL
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 18.40 0.28 ;
        RECT  17.84 -0.28 18.22 0.32 ;
        RECT  17.78 0.64 18.06 1.24 ;
        RECT  17.84 -0.28 18.00 1.24 ;
        RECT  16.74 0.64 17.02 1.24 ;
        RECT  16.80 -0.28 16.96 1.24 ;
        RECT  15.70 0.64 15.98 1.24 ;
        RECT  15.76 -0.28 15.92 1.24 ;
        RECT  14.66 0.64 14.94 1.24 ;
        RECT  14.72 -0.28 14.88 1.24 ;
        RECT  13.62 0.64 13.90 1.24 ;
        RECT  13.68 -0.28 13.84 1.24 ;
        RECT  12.62 0.88 12.90 1.16 ;
        RECT  12.68 -0.28 12.84 1.16 ;
        RECT  9.64 -0.28 9.92 0.72 ;
        RECT  5.06 -0.28 5.34 0.64 ;
        RECT  2.26 0.62 2.54 0.90 ;
        RECT  2.32 -0.28 2.48 0.90 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 18.40 3.48 ;
        RECT  17.84 2.88 18.22 3.48 ;
        RECT  17.78 1.90 18.06 2.50 ;
        RECT  17.84 1.90 18.00 3.48 ;
        RECT  16.74 1.90 17.02 2.50 ;
        RECT  16.80 1.90 16.96 3.48 ;
        RECT  15.70 1.90 15.98 2.50 ;
        RECT  15.76 1.90 15.92 3.48 ;
        RECT  14.66 1.90 14.94 2.50 ;
        RECT  14.72 1.90 14.88 3.48 ;
        RECT  13.62 1.90 13.90 2.50 ;
        RECT  13.68 1.90 13.84 3.48 ;
        RECT  12.62 1.84 12.90 2.12 ;
        RECT  12.68 1.84 12.84 3.48 ;
        RECT  11.58 1.84 11.86 2.12 ;
        RECT  11.64 1.84 11.80 3.48 ;
        RECT  10.74 1.84 10.90 3.48 ;
        RECT  10.54 1.84 10.90 2.12 ;
        RECT  5.06 2.52 5.34 3.48 ;
        RECT  3.78 2.52 4.06 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.19 0.68 0.47 0.96 ;
        RECT  0.19 1.88 0.47 2.16 ;
        RECT  0.19 0.68 0.35 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  1.67 0.62 2.02 0.90 ;
        RECT  1.53 1.12 1.83 1.40 ;
        RECT  1.67 0.62 1.83 2.20 ;
        RECT  1.67 1.92 2.02 2.20 ;
        RECT  2.78 0.62 3.10 0.90 ;
        RECT  2.94 1.22 3.22 1.50 ;
        RECT  2.94 0.62 3.10 2.20 ;
        RECT  2.78 1.92 3.10 2.20 ;
        RECT  0.71 0.68 0.99 0.96 ;
        RECT  3.26 0.76 3.54 1.04 ;
        RECT  0.77 0.68 0.93 2.16 ;
        RECT  0.71 1.88 0.99 2.16 ;
        RECT  3.38 0.76 3.54 2.26 ;
        RECT  0.83 1.88 0.99 2.52 ;
        RECT  3.26 1.98 3.42 2.52 ;
        RECT  0.83 2.36 3.42 2.52 ;
        RECT  3.90 0.44 4.90 0.60 ;
        RECT  4.62 0.44 4.90 0.72 ;
        RECT  3.90 0.44 4.06 1.04 ;
        RECT  3.74 0.76 3.90 2.26 ;
        RECT  3.74 1.98 4.06 2.26 ;
        RECT  5.82 0.96 6.26 1.24 ;
        RECT  6.10 1.46 6.42 1.74 ;
        RECT  6.10 0.96 6.26 2.20 ;
        RECT  5.82 1.92 6.26 2.20 ;
        RECT  6.42 0.44 6.70 0.72 ;
        RECT  5.50 0.56 6.70 0.72 ;
        RECT  5.50 0.56 5.66 1.12 ;
        RECT  4.82 0.96 5.66 1.12 ;
        RECT  4.82 0.96 5.10 1.24 ;
        RECT  4.90 0.96 5.06 2.20 ;
        RECT  4.78 1.92 5.06 2.20 ;
        RECT  4.78 2.04 5.66 2.20 ;
        RECT  5.50 2.04 5.66 2.64 ;
        RECT  5.50 2.48 6.70 2.64 ;
        RECT  6.42 2.48 6.70 2.76 ;
        RECT  8.02 0.88 8.30 1.16 ;
        RECT  8.02 0.88 8.18 2.12 ;
        RECT  7.80 1.84 8.18 2.12 ;
        RECT  8.50 1.84 8.78 2.12 ;
        RECT  7.80 1.96 8.78 2.12 ;
        RECT  9.20 0.44 9.48 0.72 ;
        RECT  8.66 0.56 9.48 0.72 ;
        RECT  8.54 0.88 8.82 1.16 ;
        RECT  8.66 0.56 8.82 1.68 ;
        RECT  8.66 1.52 9.10 1.68 ;
        RECT  8.94 1.52 9.10 2.12 ;
        RECT  8.94 1.84 9.30 2.12 ;
        RECT  6.98 0.87 7.26 1.15 ;
        RECT  6.42 0.99 7.26 1.15 ;
        RECT  6.42 0.96 6.70 1.24 ;
        RECT  6.58 0.99 6.74 2.12 ;
        RECT  6.55 1.84 6.83 2.12 ;
        RECT  6.55 1.96 7.12 2.12 ;
        RECT  6.96 1.96 7.12 2.76 ;
        RECT  10.30 2.42 10.58 2.76 ;
        RECT  6.96 2.60 10.58 2.76 ;
        RECT  10.50 0.50 10.78 0.78 ;
        RECT  9.06 0.88 9.34 1.20 ;
        RECT  9.68 0.92 9.96 1.20 ;
        RECT  10.50 0.50 10.66 1.20 ;
        RECT  9.06 1.04 10.66 1.20 ;
        RECT  9.46 1.04 9.62 2.12 ;
        RECT  9.46 1.84 9.82 2.12 ;
        RECT  7.48 0.87 7.78 1.15 ;
        RECT  11.16 0.92 11.44 1.20 ;
        RECT  9.98 1.52 11.32 1.68 ;
        RECT  11.16 0.92 11.32 2.12 ;
        RECT  7.36 1.84 7.64 2.12 ;
        RECT  11.06 1.84 11.34 2.12 ;
        RECT  7.48 0.87 7.64 2.44 ;
        RECT  9.98 1.52 10.14 2.44 ;
        RECT  7.48 2.28 10.14 2.44 ;
        RECT  11.72 0.88 12.00 1.16 ;
        RECT  11.72 1.00 12.27 1.16 ;
        RECT  12.11 1.46 13.10 1.62 ;
        RECT  12.82 1.40 13.10 1.68 ;
        RECT  12.11 1.00 12.27 2.12 ;
        RECT  12.10 1.84 12.38 2.12 ;
        RECT  13.14 0.88 13.42 1.16 ;
        RECT  13.14 1.84 13.42 2.12 ;
        RECT  13.26 0.88 13.42 2.76 ;
        RECT  13.17 2.48 13.45 2.76 ;
    END
END DFFDERZSP8V1_0

MACRO DFFDERZSP4V1_0
    CLASS CORE ;
    FOREIGN DFFDERZSP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.45 1.06 2.78 1.34 ;
        RECT  2.26 1.06 2.78 1.30 ;
        END
    END SEL
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.99 1.46 2.34 1.76 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 31.58  LAYER ME1  ;
        ANTENNADIFFAREA 14.14  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.18  LAYER ME1  ;
        ANTENNAMAXAREACAR 26.74  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.21 1.88 1.51 2.16 ;
        RECT  1.21 0.66 1.51 0.96 ;
        RECT  1.21 0.66 1.37 2.16 ;
        END
    END D
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 31.90  LAYER ME1  ;
        ANTENNADIFFAREA 14.14  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.18  LAYER ME1  ;
        ANTENNAMAXAREACAR 27.02  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.42 1.46 4.74 1.74 ;
        RECT  4.34 0.88 4.62 1.16 ;
        RECT  4.30 1.98 4.58 2.26 ;
        RECT  4.42 0.88 4.58 2.26 ;
        END
    END TD
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.63 1.40 5.94 1.76 ;
        END
    END CK
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.57 1.40 11.95 1.68 ;
        END
    END RB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 31.90  LAYER ME1  ;
        ANTENNADIFFAREA 14.13  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.18  LAYER ME1  ;
        ANTENNAMAXAREACAR 27.02  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.14 1.90 14.42 2.50 ;
        RECT  14.14 0.64 14.42 1.24 ;
        RECT  14.14 0.64 14.34 2.50 ;
        RECT  14.06 1.46 14.34 1.74 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 31.90  LAYER ME1  ;
        ANTENNADIFFAREA 14.38  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.18  LAYER ME1  ;
        ANTENNAMAXAREACAR 27.02  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  15.26 1.46 15.54 1.74 ;
        RECT  15.18 1.90 15.46 2.50 ;
        RECT  15.26 0.64 15.46 2.50 ;
        RECT  15.18 0.64 15.46 1.24 ;
        END
    END QB
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 16.40 3.48 ;
        RECT  15.78 2.88 16.22 3.48 ;
        RECT  15.70 1.90 15.98 2.50 ;
        RECT  15.78 1.90 15.94 3.48 ;
        RECT  14.66 1.90 14.94 2.50 ;
        RECT  14.72 1.90 14.88 3.48 ;
        RECT  13.62 1.90 13.90 2.50 ;
        RECT  13.68 1.90 13.84 3.48 ;
        RECT  12.62 1.84 12.90 2.12 ;
        RECT  12.68 1.84 12.84 3.48 ;
        RECT  11.58 1.84 11.86 2.12 ;
        RECT  11.64 1.84 11.80 3.48 ;
        RECT  10.74 1.84 10.90 3.48 ;
        RECT  10.54 1.84 10.90 2.12 ;
        RECT  5.06 2.52 5.34 3.48 ;
        RECT  3.78 2.52 4.06 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 16.40 0.28 ;
        RECT  15.78 -0.28 16.22 0.32 ;
        RECT  15.70 0.64 15.98 1.24 ;
        RECT  15.78 -0.28 15.94 1.24 ;
        RECT  14.66 0.64 14.94 1.24 ;
        RECT  14.72 -0.28 14.88 1.24 ;
        RECT  13.62 0.64 13.90 1.24 ;
        RECT  13.68 -0.28 13.84 1.24 ;
        RECT  12.62 0.88 12.90 1.16 ;
        RECT  12.68 -0.28 12.84 1.16 ;
        RECT  9.64 -0.28 9.92 0.72 ;
        RECT  5.06 -0.28 5.34 0.64 ;
        RECT  2.26 0.62 2.54 0.90 ;
        RECT  2.32 -0.28 2.48 0.90 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.19 0.68 0.47 0.96 ;
        RECT  0.19 1.88 0.47 2.16 ;
        RECT  0.19 0.68 0.35 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  1.67 0.62 2.02 0.90 ;
        RECT  1.53 1.12 1.83 1.40 ;
        RECT  1.67 0.62 1.83 2.20 ;
        RECT  1.67 1.92 2.02 2.20 ;
        RECT  2.78 0.62 3.10 0.90 ;
        RECT  2.94 1.22 3.22 1.50 ;
        RECT  2.94 0.62 3.10 2.20 ;
        RECT  2.78 1.92 3.10 2.20 ;
        RECT  0.71 0.68 0.99 0.96 ;
        RECT  3.26 0.76 3.54 1.04 ;
        RECT  0.77 0.68 0.93 2.16 ;
        RECT  0.71 1.88 0.99 2.16 ;
        RECT  3.38 0.76 3.54 2.26 ;
        RECT  0.83 1.88 0.99 2.52 ;
        RECT  3.26 1.98 3.42 2.52 ;
        RECT  0.83 2.36 3.42 2.52 ;
        RECT  3.90 0.44 4.90 0.60 ;
        RECT  4.62 0.44 4.90 0.72 ;
        RECT  3.90 0.44 4.06 1.04 ;
        RECT  3.74 0.76 3.90 2.26 ;
        RECT  3.74 1.98 4.06 2.26 ;
        RECT  5.82 0.96 6.26 1.24 ;
        RECT  6.10 1.46 6.42 1.74 ;
        RECT  6.10 0.96 6.26 2.20 ;
        RECT  5.82 1.92 6.26 2.20 ;
        RECT  6.42 0.44 6.70 0.72 ;
        RECT  5.50 0.56 6.70 0.72 ;
        RECT  5.50 0.56 5.66 1.12 ;
        RECT  4.82 0.96 5.66 1.12 ;
        RECT  4.82 0.96 5.10 1.24 ;
        RECT  4.90 0.96 5.06 2.20 ;
        RECT  4.78 1.92 5.06 2.20 ;
        RECT  4.78 2.04 5.66 2.20 ;
        RECT  5.50 2.04 5.66 2.64 ;
        RECT  5.50 2.48 6.70 2.64 ;
        RECT  6.42 2.48 6.70 2.76 ;
        RECT  8.02 0.88 8.30 1.16 ;
        RECT  8.02 0.88 8.18 2.12 ;
        RECT  7.80 1.84 8.18 2.12 ;
        RECT  8.50 1.84 8.78 2.12 ;
        RECT  7.80 1.96 8.78 2.12 ;
        RECT  9.20 0.44 9.48 0.72 ;
        RECT  8.66 0.56 9.48 0.72 ;
        RECT  8.54 0.88 8.82 1.16 ;
        RECT  8.66 0.56 8.82 1.68 ;
        RECT  8.66 1.52 9.10 1.68 ;
        RECT  8.94 1.52 9.10 2.12 ;
        RECT  8.94 1.84 9.30 2.12 ;
        RECT  6.98 0.87 7.26 1.15 ;
        RECT  6.42 0.99 7.26 1.15 ;
        RECT  6.42 0.96 6.70 1.24 ;
        RECT  6.58 0.99 6.74 2.12 ;
        RECT  6.55 1.84 6.83 2.12 ;
        RECT  6.55 1.96 7.12 2.12 ;
        RECT  6.96 1.96 7.12 2.76 ;
        RECT  10.30 2.42 10.58 2.76 ;
        RECT  6.96 2.60 10.58 2.76 ;
        RECT  10.50 0.50 10.78 0.78 ;
        RECT  9.06 0.88 9.34 1.20 ;
        RECT  9.68 0.92 9.96 1.20 ;
        RECT  10.50 0.50 10.66 1.20 ;
        RECT  9.06 1.04 10.66 1.20 ;
        RECT  9.46 1.04 9.62 2.12 ;
        RECT  9.46 1.84 9.82 2.12 ;
        RECT  7.48 0.87 7.78 1.15 ;
        RECT  11.16 0.92 11.44 1.20 ;
        RECT  9.98 1.52 11.32 1.68 ;
        RECT  11.16 0.92 11.32 2.12 ;
        RECT  7.36 1.84 7.64 2.12 ;
        RECT  11.06 1.84 11.34 2.12 ;
        RECT  7.48 0.87 7.64 2.44 ;
        RECT  9.98 1.52 10.14 2.44 ;
        RECT  7.48 2.28 10.14 2.44 ;
        RECT  11.72 0.88 12.00 1.16 ;
        RECT  11.72 1.00 12.27 1.16 ;
        RECT  12.11 1.46 13.10 1.62 ;
        RECT  12.82 1.40 13.10 1.68 ;
        RECT  12.11 1.00 12.27 2.12 ;
        RECT  12.10 1.84 12.38 2.12 ;
        RECT  13.14 0.88 13.42 1.16 ;
        RECT  13.14 1.84 13.42 2.12 ;
        RECT  13.26 0.88 13.42 2.76 ;
        RECT  13.17 2.48 13.45 2.76 ;
    END
END DFFDERZSP4V1_0

MACRO DFFDERZSP2V1_0
    CLASS CORE ;
    FOREIGN DFFDERZSP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 29.65  LAYER ME1  ;
        ANTENNADIFFAREA 12.80  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.89  LAYER ME1  ;
        ANTENNAMAXAREACAR 33.21  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.78 1.46 15.12 1.74 ;
        RECT  14.66 1.90 14.94 2.50 ;
        RECT  14.78 0.64 14.94 2.50 ;
        RECT  14.66 0.64 14.94 1.24 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 29.65  LAYER ME1  ;
        ANTENNADIFFAREA 12.80  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.89  LAYER ME1  ;
        ANTENNAMAXAREACAR 33.21  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.66 1.46 13.94 1.74 ;
        RECT  13.62 1.90 13.90 2.50 ;
        RECT  13.66 0.64 13.90 2.50 ;
        RECT  13.62 0.64 13.90 1.24 ;
        END
    END Q
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.57 1.40 11.95 1.68 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.63 1.40 5.94 1.76 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 29.65  LAYER ME1  ;
        ANTENNADIFFAREA 12.80  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.89  LAYER ME1  ;
        ANTENNAMAXAREACAR 33.21  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.42 1.46 4.74 1.74 ;
        RECT  4.34 0.88 4.62 1.16 ;
        RECT  4.30 1.98 4.58 2.26 ;
        RECT  4.42 0.88 4.58 2.26 ;
        END
    END TD
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 29.33  LAYER ME1  ;
        ANTENNADIFFAREA 12.80  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.89  LAYER ME1  ;
        ANTENNAMAXAREACAR 32.85  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.21 1.88 1.51 2.16 ;
        RECT  1.21 0.66 1.51 0.96 ;
        RECT  1.21 0.66 1.37 2.16 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.99 1.46 2.34 1.76 ;
        END
    END E
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.45 1.06 2.78 1.34 ;
        RECT  2.26 1.06 2.78 1.30 ;
        END
    END SEL
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 15.20 0.28 ;
        RECT  14.74 -0.28 15.02 0.32 ;
        RECT  14.14 0.64 14.42 1.24 ;
        RECT  14.20 -0.28 14.36 1.24 ;
        RECT  12.62 0.88 12.90 1.16 ;
        RECT  12.68 -0.28 12.84 1.16 ;
        RECT  9.64 -0.28 9.92 0.72 ;
        RECT  5.06 -0.28 5.34 0.64 ;
        RECT  2.26 0.62 2.54 0.90 ;
        RECT  2.32 -0.28 2.48 0.90 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 15.20 3.48 ;
        RECT  14.74 2.88 15.02 3.48 ;
        RECT  14.14 1.90 14.42 2.50 ;
        RECT  14.20 1.90 14.36 3.48 ;
        RECT  12.62 1.84 12.90 2.12 ;
        RECT  12.68 1.84 12.84 3.48 ;
        RECT  11.58 1.84 11.86 2.12 ;
        RECT  11.64 1.84 11.80 3.48 ;
        RECT  10.74 1.84 10.90 3.48 ;
        RECT  10.54 1.84 10.90 2.12 ;
        RECT  5.06 2.52 5.34 3.48 ;
        RECT  3.78 2.52 4.06 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.19 0.68 0.47 0.96 ;
        RECT  0.19 1.88 0.47 2.16 ;
        RECT  0.19 0.68 0.35 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  1.67 0.62 2.02 0.90 ;
        RECT  1.53 1.12 1.83 1.40 ;
        RECT  1.67 0.62 1.83 2.20 ;
        RECT  1.67 1.92 2.02 2.20 ;
        RECT  2.78 0.62 3.10 0.90 ;
        RECT  2.94 1.22 3.22 1.50 ;
        RECT  2.94 0.62 3.10 2.20 ;
        RECT  2.78 1.92 3.10 2.20 ;
        RECT  0.71 0.68 0.99 0.96 ;
        RECT  3.26 0.76 3.54 1.04 ;
        RECT  0.77 0.68 0.93 2.16 ;
        RECT  0.71 1.88 0.99 2.16 ;
        RECT  3.38 0.76 3.54 2.26 ;
        RECT  0.83 1.88 0.99 2.52 ;
        RECT  3.26 1.98 3.42 2.52 ;
        RECT  0.83 2.36 3.42 2.52 ;
        RECT  3.90 0.44 4.90 0.60 ;
        RECT  4.62 0.44 4.90 0.72 ;
        RECT  3.90 0.44 4.06 1.04 ;
        RECT  3.74 0.76 3.90 2.26 ;
        RECT  3.74 1.98 4.06 2.26 ;
        RECT  5.82 0.96 6.26 1.24 ;
        RECT  6.10 1.46 6.42 1.74 ;
        RECT  6.10 0.96 6.26 2.20 ;
        RECT  5.82 1.92 6.26 2.20 ;
        RECT  6.42 0.44 6.70 0.72 ;
        RECT  5.50 0.56 6.70 0.72 ;
        RECT  5.50 0.56 5.66 1.12 ;
        RECT  4.82 0.96 5.66 1.12 ;
        RECT  4.82 0.96 5.10 1.24 ;
        RECT  4.90 0.96 5.06 2.20 ;
        RECT  4.78 1.92 5.06 2.20 ;
        RECT  4.78 2.04 5.66 2.20 ;
        RECT  5.50 2.04 5.66 2.64 ;
        RECT  5.50 2.48 6.70 2.64 ;
        RECT  6.42 2.48 6.70 2.76 ;
        RECT  8.02 0.88 8.30 1.16 ;
        RECT  8.02 0.88 8.18 2.12 ;
        RECT  7.80 1.84 8.18 2.12 ;
        RECT  8.50 1.84 8.78 2.12 ;
        RECT  7.80 1.96 8.78 2.12 ;
        RECT  9.20 0.44 9.48 0.72 ;
        RECT  8.66 0.56 9.48 0.72 ;
        RECT  8.54 0.88 8.82 1.16 ;
        RECT  8.66 0.56 8.82 1.68 ;
        RECT  8.66 1.52 9.10 1.68 ;
        RECT  8.94 1.52 9.10 2.12 ;
        RECT  8.94 1.84 9.30 2.12 ;
        RECT  6.98 0.87 7.26 1.15 ;
        RECT  6.42 0.99 7.26 1.15 ;
        RECT  6.42 0.96 6.70 1.24 ;
        RECT  6.58 0.99 6.74 2.12 ;
        RECT  6.55 1.84 6.83 2.12 ;
        RECT  6.55 1.96 7.12 2.12 ;
        RECT  6.96 1.96 7.12 2.76 ;
        RECT  10.30 2.42 10.58 2.76 ;
        RECT  6.96 2.60 10.58 2.76 ;
        RECT  10.50 0.50 10.78 0.78 ;
        RECT  9.06 0.88 9.34 1.20 ;
        RECT  9.68 0.92 9.96 1.20 ;
        RECT  10.50 0.50 10.66 1.20 ;
        RECT  9.06 1.04 10.66 1.20 ;
        RECT  9.46 1.04 9.62 2.12 ;
        RECT  9.46 1.84 9.82 2.12 ;
        RECT  7.48 0.87 7.78 1.15 ;
        RECT  11.16 0.92 11.44 1.20 ;
        RECT  9.98 1.52 11.32 1.68 ;
        RECT  11.16 0.92 11.32 2.12 ;
        RECT  7.36 1.84 7.64 2.12 ;
        RECT  11.06 1.84 11.34 2.12 ;
        RECT  7.48 0.87 7.64 2.44 ;
        RECT  9.98 1.52 10.14 2.44 ;
        RECT  7.48 2.28 10.14 2.44 ;
        RECT  11.72 0.88 12.00 1.16 ;
        RECT  11.72 1.00 12.27 1.16 ;
        RECT  12.11 1.46 13.10 1.62 ;
        RECT  12.82 1.40 13.10 1.68 ;
        RECT  12.11 1.00 12.27 2.12 ;
        RECT  12.10 1.84 12.38 2.12 ;
        RECT  13.14 0.88 13.42 1.16 ;
        RECT  13.14 1.84 13.42 2.12 ;
        RECT  13.26 0.88 13.42 2.76 ;
        RECT  13.17 2.48 13.45 2.76 ;
    END
END DFFDERZSP2V1_0

MACRO DFFDERZSP1V1_0
    CLASS CORE ;
    FOREIGN DFFDERZSP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 28.92  LAYER ME1  ;
        ANTENNADIFFAREA 12.11  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.74  LAYER ME1  ;
        ANTENNAMAXAREACAR 39.12  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.21 1.88 1.51 2.16 ;
        RECT  1.21 0.66 1.51 0.96 ;
        RECT  1.21 0.66 1.37 2.16 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.99 1.46 2.34 1.76 ;
        END
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.63 1.40 5.94 1.76 ;
        END
    END CK
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.57 1.40 11.95 1.68 ;
        END
    END RB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 29.24  LAYER ME1  ;
        ANTENNADIFFAREA 12.11  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.74  LAYER ME1  ;
        ANTENNAMAXAREACAR 39.55  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.66 1.46 13.94 1.74 ;
        RECT  13.62 1.90 13.90 2.18 ;
        RECT  13.66 0.88 13.90 2.18 ;
        RECT  13.62 0.88 13.90 1.16 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 29.24  LAYER ME1  ;
        ANTENNADIFFAREA 12.11  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.74  LAYER ME1  ;
        ANTENNAMAXAREACAR 39.55  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.78 1.46 15.12 1.74 ;
        RECT  14.66 1.90 14.94 2.18 ;
        RECT  14.78 0.88 14.94 2.18 ;
        RECT  14.66 0.88 14.94 1.16 ;
        END
    END QB
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.45 1.06 2.78 1.34 ;
        RECT  2.26 1.06 2.78 1.30 ;
        END
    END SEL
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 29.24  LAYER ME1  ;
        ANTENNADIFFAREA 12.11  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.74  LAYER ME1  ;
        ANTENNAMAXAREACAR 39.55  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.42 1.46 4.74 1.74 ;
        RECT  4.34 0.88 4.62 1.16 ;
        RECT  4.30 1.98 4.58 2.26 ;
        RECT  4.42 0.88 4.58 2.26 ;
        END
    END TD
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 15.20 3.48 ;
        RECT  14.74 2.88 15.02 3.48 ;
        RECT  14.14 1.90 14.42 2.18 ;
        RECT  14.20 1.90 14.36 3.48 ;
        RECT  12.62 1.84 12.90 2.12 ;
        RECT  12.68 1.84 12.84 3.48 ;
        RECT  11.58 1.84 11.86 2.12 ;
        RECT  11.64 1.84 11.80 3.48 ;
        RECT  10.74 1.84 10.90 3.48 ;
        RECT  10.54 1.84 10.90 2.12 ;
        RECT  5.06 2.52 5.34 3.48 ;
        RECT  3.78 2.52 4.06 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 15.20 0.28 ;
        RECT  14.74 -0.28 15.02 0.32 ;
        RECT  14.14 0.88 14.42 1.16 ;
        RECT  14.20 -0.28 14.36 1.16 ;
        RECT  12.62 0.88 12.90 1.16 ;
        RECT  12.68 -0.28 12.84 1.16 ;
        RECT  9.64 -0.28 9.92 0.72 ;
        RECT  5.06 -0.28 5.34 0.64 ;
        RECT  2.26 0.62 2.54 0.90 ;
        RECT  2.32 -0.28 2.48 0.90 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.19 0.68 0.47 0.96 ;
        RECT  0.19 1.88 0.47 2.16 ;
        RECT  0.19 0.68 0.35 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  1.67 0.62 2.02 0.90 ;
        RECT  1.53 1.12 1.83 1.40 ;
        RECT  1.67 0.62 1.83 2.20 ;
        RECT  1.67 1.92 2.02 2.20 ;
        RECT  2.78 0.62 3.10 0.90 ;
        RECT  2.94 1.22 3.22 1.50 ;
        RECT  2.94 0.62 3.10 2.20 ;
        RECT  2.78 1.92 3.10 2.20 ;
        RECT  0.71 0.68 0.99 0.96 ;
        RECT  3.26 0.76 3.54 1.04 ;
        RECT  0.77 0.68 0.93 2.16 ;
        RECT  0.71 1.88 0.99 2.16 ;
        RECT  3.38 0.76 3.54 2.26 ;
        RECT  0.83 1.88 0.99 2.52 ;
        RECT  3.26 1.98 3.42 2.52 ;
        RECT  0.83 2.36 3.42 2.52 ;
        RECT  3.90 0.44 4.90 0.60 ;
        RECT  4.62 0.44 4.90 0.72 ;
        RECT  3.90 0.44 4.06 1.04 ;
        RECT  3.74 0.76 3.90 2.26 ;
        RECT  3.74 1.98 4.06 2.26 ;
        RECT  5.82 0.96 6.26 1.24 ;
        RECT  6.10 1.46 6.42 1.74 ;
        RECT  6.10 0.96 6.26 2.20 ;
        RECT  5.82 1.92 6.26 2.20 ;
        RECT  6.42 0.44 6.70 0.72 ;
        RECT  5.50 0.56 6.70 0.72 ;
        RECT  5.50 0.56 5.66 1.12 ;
        RECT  4.82 0.96 5.66 1.12 ;
        RECT  4.82 0.96 5.10 1.24 ;
        RECT  4.90 0.96 5.06 2.20 ;
        RECT  4.78 1.92 5.06 2.20 ;
        RECT  4.78 2.04 5.66 2.20 ;
        RECT  5.50 2.04 5.66 2.64 ;
        RECT  5.50 2.48 6.70 2.64 ;
        RECT  6.42 2.48 6.70 2.76 ;
        RECT  8.02 0.88 8.30 1.16 ;
        RECT  8.02 0.88 8.18 2.12 ;
        RECT  7.80 1.84 8.18 2.12 ;
        RECT  8.50 1.84 8.78 2.12 ;
        RECT  7.80 1.96 8.78 2.12 ;
        RECT  9.20 0.44 9.48 0.72 ;
        RECT  8.66 0.56 9.48 0.72 ;
        RECT  8.54 0.88 8.82 1.16 ;
        RECT  8.66 0.56 8.82 1.68 ;
        RECT  8.66 1.52 9.10 1.68 ;
        RECT  8.94 1.52 9.10 2.12 ;
        RECT  8.94 1.84 9.30 2.12 ;
        RECT  6.98 0.87 7.26 1.15 ;
        RECT  6.42 0.99 7.26 1.15 ;
        RECT  6.42 0.96 6.70 1.24 ;
        RECT  6.58 0.99 6.74 2.12 ;
        RECT  6.55 1.84 6.83 2.12 ;
        RECT  6.55 1.96 7.12 2.12 ;
        RECT  6.96 1.96 7.12 2.76 ;
        RECT  10.30 2.42 10.58 2.76 ;
        RECT  6.96 2.60 10.58 2.76 ;
        RECT  10.50 0.50 10.78 0.78 ;
        RECT  9.06 0.88 9.34 1.20 ;
        RECT  9.68 0.92 9.96 1.20 ;
        RECT  10.50 0.50 10.66 1.20 ;
        RECT  9.06 1.04 10.66 1.20 ;
        RECT  9.46 1.04 9.62 2.12 ;
        RECT  9.46 1.84 9.82 2.12 ;
        RECT  7.48 0.87 7.78 1.15 ;
        RECT  11.16 0.92 11.44 1.20 ;
        RECT  9.98 1.52 11.32 1.68 ;
        RECT  11.16 0.92 11.32 2.12 ;
        RECT  7.36 1.84 7.64 2.12 ;
        RECT  11.06 1.84 11.34 2.12 ;
        RECT  7.48 0.87 7.64 2.44 ;
        RECT  9.98 1.52 10.14 2.44 ;
        RECT  7.48 2.28 10.14 2.44 ;
        RECT  11.72 0.88 12.00 1.16 ;
        RECT  11.72 1.00 12.27 1.16 ;
        RECT  12.11 1.46 13.10 1.62 ;
        RECT  12.82 1.40 13.10 1.68 ;
        RECT  12.11 1.00 12.27 2.12 ;
        RECT  12.10 1.84 12.38 2.12 ;
        RECT  13.14 0.88 13.42 1.16 ;
        RECT  13.14 1.84 13.42 2.12 ;
        RECT  13.26 0.88 13.42 2.76 ;
        RECT  13.17 2.48 13.45 2.76 ;
    END
END DFFDERZSP1V1_0

MACRO DFFDERSZSP8V1_0
    CLASS CORE ;
    FOREIGN DFFDERSZSP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 20.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 38.91  LAYER ME1  ;
        ANTENNADIFFAREA 18.80  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.76  LAYER ME1  ;
        ANTENNAMAXAREACAR 22.15  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  18.90 1.90 19.18 2.50 ;
        RECT  18.90 0.64 19.18 1.24 ;
        RECT  18.90 0.64 19.06 2.50 ;
        RECT  17.98 1.52 19.06 1.68 ;
        RECT  17.98 1.46 18.34 1.74 ;
        RECT  17.86 1.90 18.14 2.50 ;
        RECT  17.98 0.64 18.14 2.50 ;
        RECT  17.86 0.64 18.14 1.24 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 38.91  LAYER ME1  ;
        ANTENNADIFFAREA 18.56  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.76  LAYER ME1  ;
        ANTENNAMAXAREACAR 22.15  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  16.82 1.90 17.10 2.50 ;
        RECT  16.82 0.64 17.10 1.24 ;
        RECT  16.82 0.64 16.98 2.50 ;
        RECT  15.66 1.52 16.98 1.68 ;
        RECT  15.78 1.90 16.06 2.50 ;
        RECT  15.78 0.64 16.06 1.24 ;
        RECT  15.78 0.64 15.94 2.50 ;
        RECT  15.66 1.46 15.94 1.74 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.06 0.44 14.34 0.94 ;
        RECT  13.80 0.44 14.34 0.72 ;
        END
    END SB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.34 1.40 12.76 1.68 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.64 1.40 5.94 1.76 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 38.59  LAYER ME1  ;
        ANTENNADIFFAREA 18.29  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.76  LAYER ME1  ;
        ANTENNAMAXAREACAR 21.97  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.21 1.88 1.51 2.16 ;
        RECT  1.21 0.66 1.51 0.96 ;
        RECT  1.21 0.66 1.37 2.16 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.99 1.46 2.34 1.76 ;
        END
    END E
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.45 1.06 2.78 1.34 ;
        RECT  2.26 1.06 2.78 1.30 ;
        END
    END SEL
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 38.91  LAYER ME1  ;
        ANTENNADIFFAREA 18.29  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.76  LAYER ME1  ;
        ANTENNAMAXAREACAR 22.15  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.42 1.46 4.74 1.74 ;
        RECT  4.42 2.42 4.72 2.70 ;
        RECT  4.34 0.88 4.62 1.16 ;
        RECT  4.42 0.88 4.58 2.70 ;
        RECT  4.30 1.98 4.58 2.26 ;
        END
    END TD
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 20.00 0.28 ;
        RECT  19.48 -0.28 19.82 0.32 ;
        RECT  19.42 0.64 19.70 1.24 ;
        RECT  19.48 -0.28 19.64 1.24 ;
        RECT  18.38 0.64 18.66 1.24 ;
        RECT  18.44 -0.28 18.60 1.24 ;
        RECT  17.34 0.64 17.62 1.24 ;
        RECT  17.40 -0.28 17.56 1.24 ;
        RECT  16.30 0.64 16.58 1.24 ;
        RECT  16.36 -0.28 16.52 1.24 ;
        RECT  15.26 0.64 15.54 1.24 ;
        RECT  15.32 -0.28 15.48 1.24 ;
        RECT  13.43 0.88 13.78 1.16 ;
        RECT  13.43 -0.28 13.59 1.16 ;
        RECT  11.04 -0.28 11.32 0.68 ;
        RECT  5.06 -0.28 5.34 0.64 ;
        RECT  2.26 0.62 2.54 0.90 ;
        RECT  2.32 -0.28 2.48 0.90 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 20.00 3.48 ;
        RECT  19.48 2.88 19.82 3.48 ;
        RECT  19.42 1.90 19.70 2.50 ;
        RECT  19.48 1.90 19.64 3.48 ;
        RECT  18.38 1.90 18.66 2.50 ;
        RECT  18.44 1.90 18.60 3.48 ;
        RECT  17.34 1.90 17.62 2.50 ;
        RECT  17.40 1.90 17.56 3.48 ;
        RECT  16.30 1.90 16.58 2.50 ;
        RECT  16.36 1.90 16.52 3.48 ;
        RECT  15.26 1.90 15.54 2.50 ;
        RECT  15.32 1.90 15.48 3.48 ;
        RECT  14.66 2.40 14.94 3.48 ;
        RECT  13.44 1.84 13.72 2.12 ;
        RECT  13.50 1.84 13.66 3.48 ;
        RECT  12.40 1.84 12.68 2.12 ;
        RECT  12.46 1.84 12.62 3.48 ;
        RECT  11.12 1.96 11.64 2.12 ;
        RECT  11.36 1.84 11.64 2.12 ;
        RECT  11.00 2.52 11.28 3.48 ;
        RECT  11.12 1.96 11.28 3.48 ;
        RECT  5.06 2.52 5.34 3.48 ;
        RECT  3.78 2.52 4.06 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.19 0.68 0.47 0.96 ;
        RECT  0.19 1.88 0.47 2.16 ;
        RECT  0.19 0.68 0.35 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  1.67 0.62 2.02 0.90 ;
        RECT  1.53 1.12 1.83 1.40 ;
        RECT  1.67 0.62 1.83 2.20 ;
        RECT  1.67 1.92 2.02 2.20 ;
        RECT  2.78 0.62 3.10 0.90 ;
        RECT  2.94 1.22 3.22 1.50 ;
        RECT  2.94 0.62 3.10 2.20 ;
        RECT  2.78 1.92 3.10 2.20 ;
        RECT  0.71 0.68 0.99 0.96 ;
        RECT  3.26 0.76 3.54 1.04 ;
        RECT  0.77 0.68 0.93 2.16 ;
        RECT  0.71 1.88 0.99 2.16 ;
        RECT  3.38 0.76 3.54 2.26 ;
        RECT  0.83 1.88 0.99 2.52 ;
        RECT  3.26 1.98 3.42 2.52 ;
        RECT  0.83 2.36 3.42 2.52 ;
        RECT  3.90 0.44 4.90 0.60 ;
        RECT  4.62 0.44 4.90 0.72 ;
        RECT  3.90 0.44 4.06 1.04 ;
        RECT  3.74 0.76 3.90 2.26 ;
        RECT  3.74 1.98 4.06 2.26 ;
        RECT  5.82 0.96 6.26 1.24 ;
        RECT  6.10 1.46 6.42 1.74 ;
        RECT  6.10 0.96 6.26 2.20 ;
        RECT  5.82 1.92 6.26 2.20 ;
        RECT  6.42 0.44 6.70 0.72 ;
        RECT  5.50 0.56 6.70 0.72 ;
        RECT  5.50 0.56 5.66 1.12 ;
        RECT  4.82 0.96 5.66 1.12 ;
        RECT  4.82 0.96 5.10 1.24 ;
        RECT  4.90 0.96 5.06 2.20 ;
        RECT  4.78 1.92 5.06 2.20 ;
        RECT  4.78 2.04 5.66 2.20 ;
        RECT  5.50 2.04 5.66 2.64 ;
        RECT  5.50 2.48 6.60 2.64 ;
        RECT  6.32 2.48 6.60 2.76 ;
        RECT  7.94 0.88 8.26 1.16 ;
        RECT  7.94 0.88 8.10 2.00 ;
        RECT  7.60 1.84 8.58 2.00 ;
        RECT  7.60 1.84 7.88 2.12 ;
        RECT  8.30 1.84 8.58 2.12 ;
        RECT  8.50 0.88 8.78 1.16 ;
        RECT  8.62 0.88 8.78 1.58 ;
        RECT  9.46 1.14 9.74 1.58 ;
        RECT  8.62 1.42 9.74 1.58 ;
        RECT  8.74 1.42 8.90 2.12 ;
        RECT  8.74 1.84 9.10 2.12 ;
        RECT  7.10 0.50 10.50 0.66 ;
        RECT  10.22 0.50 10.50 0.78 ;
        RECT  6.98 0.86 7.26 1.14 ;
        RECT  7.10 0.50 7.26 1.14 ;
        RECT  6.42 0.98 7.26 1.14 ;
        RECT  6.42 0.96 6.70 1.24 ;
        RECT  6.64 0.98 6.80 2.12 ;
        RECT  6.64 1.84 6.92 2.12 ;
        RECT  11.48 0.50 11.76 0.78 ;
        RECT  9.02 0.82 10.06 0.98 ;
        RECT  9.02 0.82 9.30 1.16 ;
        RECT  11.48 0.50 11.64 1.16 ;
        RECT  9.90 1.00 11.64 1.16 ;
        RECT  9.90 0.96 10.26 1.24 ;
        RECT  10.20 1.00 10.36 2.12 ;
        RECT  9.34 1.84 9.62 2.12 ;
        RECT  10.20 1.84 10.54 2.12 ;
        RECT  9.34 1.96 10.54 2.12 ;
        RECT  7.42 0.86 7.78 1.14 ;
        RECT  12.02 0.96 12.46 1.24 ;
        RECT  7.42 0.86 7.58 1.48 ;
        RECT  10.70 1.52 12.18 1.68 ;
        RECT  7.16 1.84 7.44 2.12 ;
        RECT  12.02 0.96 12.18 2.12 ;
        RECT  11.88 1.84 12.18 2.12 ;
        RECT  7.28 1.32 7.44 2.44 ;
        RECT  10.70 1.52 10.86 2.44 ;
        RECT  7.28 2.28 10.86 2.44 ;
        RECT  12.66 0.88 13.08 1.16 ;
        RECT  12.92 1.46 14.46 1.62 ;
        RECT  14.18 1.40 14.46 1.68 ;
        RECT  12.92 0.88 13.08 2.12 ;
        RECT  12.92 1.84 13.20 2.12 ;
        RECT  14.50 0.88 14.82 1.16 ;
        RECT  14.66 0.88 14.82 2.16 ;
        RECT  14.66 1.88 14.94 2.16 ;
        RECT  14.17 2.00 14.94 2.16 ;
        RECT  14.17 2.00 14.33 2.76 ;
        RECT  14.05 2.48 14.33 2.76 ;
    END
END DFFDERSZSP8V1_0

MACRO DFFDERSZSP4V1_0
    CLASS CORE ;
    FOREIGN DFFDERSZSP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 34.65  LAYER ME1  ;
        ANTENNADIFFAREA 15.73  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.18  LAYER ME1  ;
        ANTENNAMAXAREACAR 29.35  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.42 1.46 4.74 1.74 ;
        RECT  4.42 2.42 4.72 2.70 ;
        RECT  4.34 0.88 4.62 1.16 ;
        RECT  4.42 0.88 4.58 2.70 ;
        RECT  4.30 1.98 4.58 2.26 ;
        END
    END TD
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.45 1.06 2.78 1.34 ;
        RECT  2.26 1.06 2.78 1.30 ;
        END
    END SEL
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.99 1.46 2.34 1.76 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 34.33  LAYER ME1  ;
        ANTENNADIFFAREA 15.73  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.18  LAYER ME1  ;
        ANTENNAMAXAREACAR 29.08  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.21 1.88 1.51 2.16 ;
        RECT  1.21 0.66 1.51 0.96 ;
        RECT  1.21 0.66 1.37 2.16 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.64 1.40 5.94 1.76 ;
        END
    END CK
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.34 1.40 12.76 1.68 ;
        END
    END RB
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.06 0.44 14.34 0.94 ;
        RECT  13.80 0.44 14.34 0.72 ;
        END
    END SB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 34.65  LAYER ME1  ;
        ANTENNADIFFAREA 15.52  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.18  LAYER ME1  ;
        ANTENNAMAXAREACAR 29.35  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  15.78 1.89 16.06 2.49 ;
        RECT  15.78 0.64 16.06 1.24 ;
        RECT  15.78 0.64 15.94 2.49 ;
        RECT  15.66 1.46 15.94 1.74 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 34.65  LAYER ME1  ;
        ANTENNADIFFAREA 15.76  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.18  LAYER ME1  ;
        ANTENNAMAXAREACAR 29.35  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  16.86 1.46 17.14 1.74 ;
        RECT  16.82 1.89 17.10 2.49 ;
        RECT  16.86 0.64 17.10 2.49 ;
        RECT  16.82 0.64 17.10 1.24 ;
        END
    END QB
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 18.00 3.48 ;
        RECT  17.40 2.88 17.82 3.48 ;
        RECT  17.34 1.89 17.62 2.49 ;
        RECT  17.40 1.89 17.56 3.48 ;
        RECT  16.30 1.89 16.58 2.49 ;
        RECT  16.36 1.89 16.52 3.48 ;
        RECT  15.26 1.89 15.54 2.49 ;
        RECT  15.32 1.89 15.48 3.48 ;
        RECT  14.66 2.40 14.94 3.48 ;
        RECT  13.44 1.84 13.72 2.12 ;
        RECT  13.50 1.84 13.66 3.48 ;
        RECT  12.40 1.84 12.68 2.12 ;
        RECT  12.46 1.84 12.62 3.48 ;
        RECT  11.12 1.96 11.64 2.12 ;
        RECT  11.36 1.84 11.64 2.12 ;
        RECT  11.00 2.52 11.28 3.48 ;
        RECT  11.12 1.96 11.28 3.48 ;
        RECT  5.06 2.52 5.34 3.48 ;
        RECT  3.78 2.52 4.06 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 18.00 0.28 ;
        RECT  17.40 -0.28 17.82 0.32 ;
        RECT  17.34 0.64 17.62 1.24 ;
        RECT  17.40 -0.28 17.56 1.24 ;
        RECT  16.30 0.64 16.58 1.24 ;
        RECT  16.36 -0.28 16.52 1.24 ;
        RECT  15.26 0.64 15.54 1.24 ;
        RECT  15.32 -0.28 15.48 1.24 ;
        RECT  13.43 0.88 13.78 1.16 ;
        RECT  13.43 -0.28 13.59 1.16 ;
        RECT  11.04 -0.28 11.32 0.68 ;
        RECT  5.06 -0.28 5.34 0.64 ;
        RECT  2.26 0.62 2.54 0.90 ;
        RECT  2.32 -0.28 2.48 0.90 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.19 0.68 0.47 0.96 ;
        RECT  0.19 1.88 0.47 2.16 ;
        RECT  0.19 0.68 0.35 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  1.67 0.62 2.02 0.90 ;
        RECT  1.53 1.12 1.83 1.40 ;
        RECT  1.67 0.62 1.83 2.20 ;
        RECT  1.67 1.92 2.02 2.20 ;
        RECT  2.78 0.62 3.10 0.90 ;
        RECT  2.94 1.22 3.22 1.50 ;
        RECT  2.94 0.62 3.10 2.20 ;
        RECT  2.78 1.92 3.10 2.20 ;
        RECT  0.71 0.68 0.99 0.96 ;
        RECT  3.26 0.76 3.54 1.04 ;
        RECT  0.77 0.68 0.93 2.16 ;
        RECT  0.71 1.88 0.99 2.16 ;
        RECT  3.38 0.76 3.54 2.26 ;
        RECT  0.83 1.88 0.99 2.52 ;
        RECT  3.26 1.98 3.42 2.52 ;
        RECT  0.83 2.36 3.42 2.52 ;
        RECT  3.90 0.44 4.90 0.60 ;
        RECT  4.62 0.44 4.90 0.72 ;
        RECT  3.90 0.44 4.06 1.04 ;
        RECT  3.74 0.76 3.90 2.26 ;
        RECT  3.74 1.98 4.06 2.26 ;
        RECT  5.82 0.96 6.26 1.24 ;
        RECT  6.10 1.46 6.42 1.74 ;
        RECT  6.10 0.96 6.26 2.20 ;
        RECT  5.82 1.92 6.26 2.20 ;
        RECT  6.42 0.44 6.70 0.72 ;
        RECT  5.50 0.56 6.70 0.72 ;
        RECT  5.50 0.56 5.66 1.12 ;
        RECT  4.82 0.96 5.66 1.12 ;
        RECT  4.82 0.96 5.10 1.24 ;
        RECT  4.90 0.96 5.06 2.20 ;
        RECT  4.78 1.92 5.06 2.20 ;
        RECT  4.78 2.04 5.66 2.20 ;
        RECT  5.50 2.04 5.66 2.64 ;
        RECT  5.50 2.48 6.60 2.64 ;
        RECT  6.32 2.48 6.60 2.76 ;
        RECT  7.94 0.88 8.26 1.16 ;
        RECT  7.94 0.88 8.10 2.00 ;
        RECT  7.60 1.84 8.58 2.00 ;
        RECT  7.60 1.84 7.88 2.12 ;
        RECT  8.30 1.84 8.58 2.12 ;
        RECT  8.50 0.88 8.78 1.16 ;
        RECT  8.62 0.88 8.78 1.58 ;
        RECT  9.46 1.14 9.74 1.58 ;
        RECT  8.62 1.42 9.74 1.58 ;
        RECT  8.74 1.42 8.90 2.12 ;
        RECT  8.74 1.84 9.10 2.12 ;
        RECT  7.10 0.50 10.50 0.66 ;
        RECT  10.22 0.50 10.50 0.78 ;
        RECT  6.98 0.86 7.26 1.14 ;
        RECT  7.10 0.50 7.26 1.14 ;
        RECT  6.42 0.98 7.26 1.14 ;
        RECT  6.42 0.96 6.70 1.24 ;
        RECT  6.64 0.98 6.80 2.12 ;
        RECT  6.64 1.84 6.92 2.12 ;
        RECT  11.48 0.50 11.76 0.78 ;
        RECT  9.02 0.82 10.06 0.98 ;
        RECT  9.02 0.82 9.30 1.16 ;
        RECT  11.48 0.50 11.64 1.16 ;
        RECT  9.90 1.00 11.64 1.16 ;
        RECT  9.90 0.96 10.26 1.24 ;
        RECT  10.20 1.00 10.36 2.12 ;
        RECT  9.34 1.84 9.62 2.12 ;
        RECT  10.20 1.84 10.54 2.12 ;
        RECT  9.34 1.96 10.54 2.12 ;
        RECT  7.42 0.86 7.78 1.14 ;
        RECT  12.02 0.96 12.46 1.24 ;
        RECT  7.42 0.86 7.58 1.48 ;
        RECT  10.70 1.52 12.18 1.68 ;
        RECT  7.16 1.84 7.44 2.12 ;
        RECT  12.02 0.96 12.18 2.12 ;
        RECT  11.88 1.84 12.18 2.12 ;
        RECT  7.28 1.32 7.44 2.44 ;
        RECT  10.70 1.52 10.86 2.44 ;
        RECT  7.28 2.28 10.86 2.44 ;
        RECT  12.66 0.88 13.08 1.16 ;
        RECT  12.92 1.46 14.46 1.62 ;
        RECT  14.18 1.40 14.46 1.68 ;
        RECT  12.92 0.88 13.08 2.12 ;
        RECT  12.92 1.84 13.20 2.12 ;
        RECT  14.50 0.88 14.82 1.16 ;
        RECT  14.66 0.88 14.82 2.16 ;
        RECT  14.66 1.88 14.94 2.16 ;
        RECT  14.17 2.00 14.94 2.16 ;
        RECT  14.17 2.00 14.33 2.76 ;
        RECT  14.05 2.48 14.33 2.76 ;
    END
END DFFDERSZSP4V1_0

MACRO DFFDERSZSP2V1_0
    CLASS CORE ;
    FOREIGN DFFDERSZSP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 32.09  LAYER ME1  ;
        ANTENNADIFFAREA 14.39  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.89  LAYER ME1  ;
        ANTENNAMAXAREACAR 35.94  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.21 1.88 1.51 2.16 ;
        RECT  1.21 0.66 1.51 0.96 ;
        RECT  1.21 0.66 1.37 2.16 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.99 1.46 2.34 1.76 ;
        END
    END E
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 32.41  LAYER ME1  ;
        ANTENNADIFFAREA 14.18  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.89  LAYER ME1  ;
        ANTENNAMAXAREACAR 36.30  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  16.42 1.46 16.72 1.74 ;
        RECT  16.30 1.89 16.58 2.49 ;
        RECT  16.42 0.64 16.58 2.49 ;
        RECT  16.30 0.64 16.58 1.24 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 32.41  LAYER ME1  ;
        ANTENNADIFFAREA 14.18  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.89  LAYER ME1  ;
        ANTENNAMAXAREACAR 36.30  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  15.26 0.64 15.54 2.49 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.06 0.44 14.34 0.94 ;
        RECT  13.80 0.44 14.34 0.72 ;
        END
    END SB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.34 1.40 12.76 1.68 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.64 1.40 5.94 1.76 ;
        END
    END CK
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.45 1.06 2.78 1.34 ;
        RECT  2.26 1.06 2.78 1.30 ;
        END
    END SEL
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 32.41  LAYER ME1  ;
        ANTENNADIFFAREA 14.39  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.89  LAYER ME1  ;
        ANTENNAMAXAREACAR 36.30  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.42 1.46 4.74 1.74 ;
        RECT  4.42 2.42 4.72 2.70 ;
        RECT  4.34 0.88 4.62 1.16 ;
        RECT  4.42 0.88 4.58 2.70 ;
        RECT  4.30 1.98 4.58 2.26 ;
        END
    END TD
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 16.80 0.28 ;
        RECT  16.34 -0.28 16.62 0.32 ;
        RECT  15.78 0.64 16.06 1.24 ;
        RECT  15.84 -0.28 16.00 1.24 ;
        RECT  13.43 0.88 13.78 1.16 ;
        RECT  13.43 -0.28 13.59 1.16 ;
        RECT  11.04 -0.28 11.32 0.68 ;
        RECT  5.06 -0.28 5.34 0.64 ;
        RECT  2.26 0.62 2.54 0.90 ;
        RECT  2.32 -0.28 2.48 0.90 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 16.80 3.48 ;
        RECT  16.34 2.88 16.62 3.48 ;
        RECT  15.78 1.89 16.06 2.49 ;
        RECT  15.84 1.89 16.00 3.48 ;
        RECT  14.66 2.40 14.94 3.48 ;
        RECT  13.44 1.84 13.72 2.12 ;
        RECT  13.50 1.84 13.66 3.48 ;
        RECT  12.40 1.84 12.68 2.12 ;
        RECT  12.46 1.84 12.62 3.48 ;
        RECT  11.12 1.96 11.64 2.12 ;
        RECT  11.36 1.84 11.64 2.12 ;
        RECT  11.00 2.52 11.28 3.48 ;
        RECT  11.12 1.96 11.28 3.48 ;
        RECT  5.06 2.52 5.34 3.48 ;
        RECT  3.78 2.52 4.06 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.19 0.68 0.47 0.96 ;
        RECT  0.19 1.88 0.47 2.16 ;
        RECT  0.19 0.68 0.35 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  1.67 0.62 2.02 0.90 ;
        RECT  1.53 1.12 1.83 1.40 ;
        RECT  1.67 0.62 1.83 2.20 ;
        RECT  1.67 1.92 2.02 2.20 ;
        RECT  2.78 0.62 3.10 0.90 ;
        RECT  2.94 1.22 3.22 1.50 ;
        RECT  2.94 0.62 3.10 2.20 ;
        RECT  2.78 1.92 3.10 2.20 ;
        RECT  0.71 0.68 0.99 0.96 ;
        RECT  3.26 0.76 3.54 1.04 ;
        RECT  0.77 0.68 0.93 2.16 ;
        RECT  0.71 1.88 0.99 2.16 ;
        RECT  3.38 0.76 3.54 2.26 ;
        RECT  0.83 1.88 0.99 2.52 ;
        RECT  3.26 1.98 3.42 2.52 ;
        RECT  0.83 2.36 3.42 2.52 ;
        RECT  3.90 0.44 4.90 0.60 ;
        RECT  4.62 0.44 4.90 0.72 ;
        RECT  3.90 0.44 4.06 1.04 ;
        RECT  3.74 0.76 3.90 2.26 ;
        RECT  3.74 1.98 4.06 2.26 ;
        RECT  5.82 0.96 6.26 1.24 ;
        RECT  6.10 1.46 6.42 1.74 ;
        RECT  6.10 0.96 6.26 2.20 ;
        RECT  5.82 1.92 6.26 2.20 ;
        RECT  6.42 0.44 6.70 0.72 ;
        RECT  5.50 0.56 6.70 0.72 ;
        RECT  5.50 0.56 5.66 1.12 ;
        RECT  4.82 0.96 5.66 1.12 ;
        RECT  4.82 0.96 5.10 1.24 ;
        RECT  4.90 0.96 5.06 2.20 ;
        RECT  4.78 1.92 5.06 2.20 ;
        RECT  4.78 2.04 5.66 2.20 ;
        RECT  5.50 2.04 5.66 2.64 ;
        RECT  5.50 2.48 6.60 2.64 ;
        RECT  6.32 2.48 6.60 2.76 ;
        RECT  7.94 0.88 8.26 1.16 ;
        RECT  7.94 0.88 8.10 2.00 ;
        RECT  7.60 1.84 8.58 2.00 ;
        RECT  7.60 1.84 7.88 2.12 ;
        RECT  8.30 1.84 8.58 2.12 ;
        RECT  8.50 0.88 8.78 1.16 ;
        RECT  8.62 0.88 8.78 1.58 ;
        RECT  9.46 1.14 9.74 1.58 ;
        RECT  8.62 1.42 9.74 1.58 ;
        RECT  8.74 1.42 8.90 2.12 ;
        RECT  8.74 1.84 9.10 2.12 ;
        RECT  7.10 0.50 10.50 0.66 ;
        RECT  10.22 0.50 10.50 0.78 ;
        RECT  6.98 0.86 7.26 1.14 ;
        RECT  7.10 0.50 7.26 1.14 ;
        RECT  6.42 0.98 7.26 1.14 ;
        RECT  6.42 0.96 6.70 1.24 ;
        RECT  6.64 0.98 6.80 2.12 ;
        RECT  6.64 1.84 6.92 2.12 ;
        RECT  11.48 0.50 11.76 0.78 ;
        RECT  9.02 0.82 10.06 0.98 ;
        RECT  9.02 0.82 9.30 1.16 ;
        RECT  11.48 0.50 11.64 1.16 ;
        RECT  9.90 1.00 11.64 1.16 ;
        RECT  9.90 0.96 10.26 1.24 ;
        RECT  10.20 1.00 10.36 2.12 ;
        RECT  9.34 1.84 9.62 2.12 ;
        RECT  10.20 1.84 10.54 2.12 ;
        RECT  9.34 1.96 10.54 2.12 ;
        RECT  7.42 0.86 7.78 1.14 ;
        RECT  12.02 0.96 12.46 1.24 ;
        RECT  7.42 0.86 7.58 1.48 ;
        RECT  10.70 1.52 12.18 1.68 ;
        RECT  7.16 1.84 7.44 2.12 ;
        RECT  12.02 0.96 12.18 2.12 ;
        RECT  11.88 1.84 12.18 2.12 ;
        RECT  7.28 1.32 7.44 2.44 ;
        RECT  10.70 1.52 10.86 2.44 ;
        RECT  7.28 2.28 10.86 2.44 ;
        RECT  12.66 0.88 13.08 1.16 ;
        RECT  12.92 1.46 14.46 1.62 ;
        RECT  14.18 1.40 14.46 1.68 ;
        RECT  12.92 0.88 13.08 2.12 ;
        RECT  12.92 1.84 13.20 2.12 ;
        RECT  14.50 0.88 14.82 1.16 ;
        RECT  14.66 0.88 14.82 2.16 ;
        RECT  14.66 1.88 14.94 2.16 ;
        RECT  14.17 2.00 14.94 2.16 ;
        RECT  14.17 2.00 14.33 2.76 ;
        RECT  14.05 2.48 14.33 2.76 ;
    END
END DFFDERSZSP2V1_0

MACRO DFFDERSZSP1V1_0
    CLASS CORE ;
    FOREIGN DFFDERSZSP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 31.86  LAYER ME1  ;
        ANTENNADIFFAREA 13.42  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.74  LAYER ME1  ;
        ANTENNAMAXAREACAR 43.10  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  16.12 1.89 16.40 2.17 ;
        RECT  16.12 0.88 16.40 1.16 ;
        RECT  16.12 0.88 16.34 2.17 ;
        RECT  16.06 1.46 16.34 1.74 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 31.86  LAYER ME1  ;
        ANTENNADIFFAREA 13.42  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.74  LAYER ME1  ;
        ANTENNAMAXAREACAR 43.10  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  15.20 1.46 15.54 1.74 ;
        RECT  15.08 1.89 15.36 2.17 ;
        RECT  15.20 0.88 15.36 2.17 ;
        RECT  15.08 0.88 15.36 1.16 ;
        END
    END Q
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.34 1.40 12.76 1.68 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.64 1.40 5.94 1.76 ;
        END
    END CK
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.06 0.44 14.34 0.94 ;
        RECT  13.80 0.44 14.34 0.72 ;
        END
    END SB
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 31.54  LAYER ME1  ;
        ANTENNADIFFAREA 13.62  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.74  LAYER ME1  ;
        ANTENNAMAXAREACAR 42.66  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.21 1.88 1.51 2.16 ;
        RECT  1.21 0.66 1.51 0.96 ;
        RECT  1.21 0.66 1.37 2.16 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.99 1.46 2.34 1.76 ;
        END
    END E
    PIN TD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 31.86  LAYER ME1  ;
        ANTENNADIFFAREA 13.62  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.74  LAYER ME1  ;
        ANTENNAMAXAREACAR 43.10  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.42 1.46 4.74 1.74 ;
        RECT  4.34 0.88 4.62 1.16 ;
        RECT  4.30 1.98 4.58 2.26 ;
        RECT  4.42 0.88 4.58 2.26 ;
        END
    END TD
    PIN SEL
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.45 1.06 2.78 1.34 ;
        RECT  2.26 1.06 2.78 1.30 ;
        END
    END SEL
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 16.80 3.48 ;
        RECT  16.34 2.88 16.62 3.48 ;
        RECT  15.60 1.89 15.88 2.17 ;
        RECT  15.66 1.89 15.82 3.48 ;
        RECT  14.28 2.52 14.56 3.48 ;
        RECT  13.44 1.84 13.72 2.12 ;
        RECT  13.50 1.84 13.66 3.48 ;
        RECT  12.40 1.84 12.68 2.12 ;
        RECT  12.46 1.84 12.62 3.48 ;
        RECT  11.12 1.96 11.64 2.12 ;
        RECT  11.36 1.84 11.64 2.12 ;
        RECT  11.00 2.52 11.28 3.48 ;
        RECT  11.12 1.96 11.28 3.48 ;
        RECT  5.06 2.52 5.34 3.48 ;
        RECT  3.78 2.52 4.06 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 16.80 0.28 ;
        RECT  16.34 -0.28 16.62 0.32 ;
        RECT  15.60 0.88 15.88 1.16 ;
        RECT  15.66 -0.28 15.82 1.16 ;
        RECT  13.43 0.88 13.78 1.16 ;
        RECT  13.43 -0.28 13.59 1.16 ;
        RECT  11.04 -0.28 11.32 0.68 ;
        RECT  5.06 -0.28 5.34 0.64 ;
        RECT  2.26 0.62 2.54 0.90 ;
        RECT  2.32 -0.28 2.48 0.90 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.19 0.68 0.47 0.96 ;
        RECT  0.19 1.88 0.47 2.16 ;
        RECT  0.19 0.68 0.35 2.76 ;
        RECT  0.10 2.48 0.38 2.76 ;
        RECT  1.67 0.62 2.02 0.90 ;
        RECT  1.53 1.12 1.83 1.40 ;
        RECT  1.67 0.62 1.83 2.20 ;
        RECT  1.67 1.92 2.02 2.20 ;
        RECT  2.78 0.62 3.10 0.90 ;
        RECT  2.94 1.22 3.22 1.50 ;
        RECT  2.94 0.62 3.10 2.20 ;
        RECT  2.78 1.92 3.10 2.20 ;
        RECT  0.71 0.68 0.99 0.96 ;
        RECT  3.26 0.76 3.54 1.04 ;
        RECT  0.77 0.68 0.93 2.16 ;
        RECT  0.71 1.88 0.99 2.16 ;
        RECT  3.38 0.76 3.54 2.26 ;
        RECT  0.83 1.88 0.99 2.52 ;
        RECT  3.26 1.98 3.42 2.52 ;
        RECT  0.83 2.36 3.42 2.52 ;
        RECT  3.90 0.44 4.90 0.60 ;
        RECT  4.62 0.44 4.90 0.72 ;
        RECT  3.90 0.44 4.06 1.04 ;
        RECT  3.74 0.76 3.90 2.26 ;
        RECT  3.74 1.98 4.06 2.26 ;
        RECT  5.82 0.96 6.26 1.24 ;
        RECT  6.10 1.46 6.42 1.74 ;
        RECT  6.10 0.96 6.26 2.20 ;
        RECT  5.82 1.92 6.26 2.20 ;
        RECT  6.42 0.44 6.70 0.72 ;
        RECT  5.50 0.56 6.70 0.72 ;
        RECT  5.50 0.56 5.66 1.12 ;
        RECT  4.82 0.96 5.66 1.12 ;
        RECT  4.82 0.96 5.10 1.24 ;
        RECT  4.90 0.96 5.06 2.20 ;
        RECT  4.78 1.92 5.06 2.20 ;
        RECT  4.78 2.04 5.66 2.20 ;
        RECT  5.50 2.04 5.66 2.64 ;
        RECT  5.50 2.48 6.60 2.64 ;
        RECT  6.32 2.48 6.60 2.76 ;
        RECT  7.94 0.88 8.26 1.16 ;
        RECT  7.94 0.88 8.10 2.00 ;
        RECT  7.60 1.84 8.58 2.00 ;
        RECT  7.60 1.84 7.88 2.12 ;
        RECT  8.30 1.84 8.58 2.12 ;
        RECT  8.50 0.88 8.78 1.16 ;
        RECT  8.62 0.88 8.78 1.58 ;
        RECT  9.46 1.14 9.74 1.58 ;
        RECT  8.62 1.42 9.74 1.58 ;
        RECT  8.74 1.42 8.90 2.12 ;
        RECT  8.74 1.84 9.10 2.12 ;
        RECT  7.10 0.50 10.50 0.66 ;
        RECT  10.22 0.50 10.50 0.78 ;
        RECT  6.98 0.86 7.26 1.14 ;
        RECT  7.10 0.50 7.26 1.14 ;
        RECT  6.42 0.98 7.26 1.14 ;
        RECT  6.42 0.96 6.70 1.24 ;
        RECT  6.64 0.98 6.80 2.12 ;
        RECT  6.64 1.84 6.92 2.12 ;
        RECT  11.48 0.50 11.76 0.78 ;
        RECT  9.02 0.82 10.06 0.98 ;
        RECT  9.02 0.82 9.30 1.16 ;
        RECT  11.48 0.50 11.64 1.16 ;
        RECT  9.90 1.00 11.64 1.16 ;
        RECT  9.90 0.96 10.26 1.24 ;
        RECT  10.20 1.00 10.36 2.12 ;
        RECT  9.34 1.84 9.62 2.12 ;
        RECT  10.20 1.84 10.54 2.12 ;
        RECT  9.34 1.96 10.54 2.12 ;
        RECT  7.42 0.86 7.78 1.14 ;
        RECT  12.02 0.96 12.46 1.24 ;
        RECT  7.42 0.86 7.58 1.48 ;
        RECT  10.70 1.52 12.18 1.68 ;
        RECT  7.16 1.84 7.44 2.12 ;
        RECT  12.02 0.96 12.18 2.12 ;
        RECT  11.88 1.84 12.18 2.12 ;
        RECT  7.28 1.32 7.44 2.44 ;
        RECT  10.70 1.52 10.86 2.44 ;
        RECT  7.28 2.28 10.86 2.44 ;
        RECT  12.66 0.88 13.08 1.16 ;
        RECT  12.92 1.46 14.46 1.62 ;
        RECT  14.18 1.40 14.46 1.68 ;
        RECT  12.92 0.88 13.08 2.12 ;
        RECT  12.92 1.84 13.20 2.12 ;
        RECT  14.50 0.88 14.78 1.16 ;
        RECT  14.62 0.88 14.78 2.16 ;
        RECT  14.28 2.00 14.88 2.16 ;
        RECT  14.28 2.00 14.56 2.28 ;
        RECT  14.72 2.00 14.88 2.64 ;
        RECT  14.72 2.48 15.26 2.64 ;
        RECT  14.98 2.48 15.26 2.76 ;
    END
END DFFDERSZSP1V1_0

MACRO DFFDERSSP8V1_0
    CLASS CORE ;
    FOREIGN DFFDERSSP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 17.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 34.20  LAYER ME1  ;
        ANTENNADIFFAREA 16.80  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.69  LAYER ME1  ;
        ANTENNAMAXAREACAR 20.24  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  16.55 1.90 16.83 2.50 ;
        RECT  16.55 0.64 16.83 1.24 ;
        RECT  16.55 0.64 16.71 2.50 ;
        RECT  15.63 1.52 16.71 1.68 ;
        RECT  15.63 1.46 15.95 1.74 ;
        RECT  15.51 1.90 15.79 2.50 ;
        RECT  15.63 0.64 15.79 2.50 ;
        RECT  15.51 0.64 15.79 1.24 ;
        END
    END QB
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 33.84  LAYER ME1  ;
        ANTENNADIFFAREA 16.28  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.69  LAYER ME1  ;
        ANTENNAMAXAREACAR 20.03  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.88 1.19 2.32 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 2.04 1.19 2.32 ;
        RECT  0.91 0.88 1.19 1.16 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.24 1.40 3.54 1.76 ;
        END
    END CK
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.99 1.40 10.41 1.68 ;
        END
    END RB
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.66 0.44 11.94 0.94 ;
        RECT  11.45 0.44 11.94 0.72 ;
        END
    END SB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 34.20  LAYER ME1  ;
        ANTENNADIFFAREA 16.56  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.69  LAYER ME1  ;
        ANTENNAMAXAREACAR 20.24  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.47 1.90 14.75 2.50 ;
        RECT  14.47 0.64 14.75 1.24 ;
        RECT  14.47 0.64 14.63 2.50 ;
        RECT  13.55 1.52 14.63 1.68 ;
        RECT  13.55 1.46 13.94 1.74 ;
        RECT  13.43 1.90 13.71 2.50 ;
        RECT  13.55 0.64 13.71 2.50 ;
        RECT  13.43 0.64 13.71 1.24 ;
        END
    END Q
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 17.60 3.48 ;
        RECT  17.13 2.88 17.42 3.48 ;
        RECT  17.07 1.90 17.35 2.50 ;
        RECT  17.13 1.90 17.29 3.48 ;
        RECT  16.03 1.90 16.31 2.50 ;
        RECT  16.09 1.90 16.25 3.48 ;
        RECT  14.99 1.90 15.27 2.50 ;
        RECT  15.05 1.90 15.21 3.48 ;
        RECT  13.95 1.90 14.23 2.50 ;
        RECT  14.01 1.90 14.17 3.48 ;
        RECT  12.91 1.90 13.19 2.50 ;
        RECT  12.97 1.90 13.13 3.48 ;
        RECT  12.31 2.40 12.59 3.48 ;
        RECT  11.09 1.84 11.37 2.12 ;
        RECT  11.15 1.84 11.31 3.48 ;
        RECT  10.05 1.84 10.33 2.12 ;
        RECT  10.11 1.84 10.27 3.48 ;
        RECT  8.77 1.96 9.29 2.12 ;
        RECT  9.01 1.84 9.29 2.12 ;
        RECT  8.65 2.52 8.93 3.48 ;
        RECT  8.77 1.96 8.93 3.48 ;
        RECT  2.71 2.52 2.99 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 17.60 0.28 ;
        RECT  17.13 -0.28 17.42 0.32 ;
        RECT  17.07 0.64 17.35 1.24 ;
        RECT  17.13 -0.28 17.29 1.24 ;
        RECT  16.03 0.64 16.31 1.24 ;
        RECT  16.09 -0.28 16.25 1.24 ;
        RECT  14.99 0.64 15.27 1.24 ;
        RECT  15.05 -0.28 15.21 1.24 ;
        RECT  13.95 0.64 14.23 1.24 ;
        RECT  14.01 -0.28 14.17 1.24 ;
        RECT  12.91 0.64 13.19 1.24 ;
        RECT  12.97 -0.28 13.13 1.24 ;
        RECT  11.08 0.88 11.43 1.16 ;
        RECT  11.08 -0.28 11.24 1.16 ;
        RECT  8.69 -0.28 8.97 0.68 ;
        RECT  2.71 -0.28 2.99 0.64 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.95 0.88 2.23 1.16 ;
        RECT  1.95 2.04 2.23 2.32 ;
        RECT  2.07 0.88 2.23 2.70 ;
        RECT  2.07 2.42 2.37 2.70 ;
        RECT  2.27 0.44 2.55 0.72 ;
        RECT  1.55 0.56 2.55 0.72 ;
        RECT  1.55 0.56 1.71 1.16 ;
        RECT  1.43 0.88 1.71 1.16 ;
        RECT  1.49 0.88 1.65 2.32 ;
        RECT  1.43 2.04 1.71 2.32 ;
        RECT  3.47 0.96 3.86 1.24 ;
        RECT  3.70 1.46 4.02 1.74 ;
        RECT  3.70 0.96 3.86 2.20 ;
        RECT  3.47 1.92 3.86 2.20 ;
        RECT  4.07 0.44 4.35 0.72 ;
        RECT  3.15 0.56 4.35 0.72 ;
        RECT  3.15 0.56 3.31 1.12 ;
        RECT  2.43 0.96 3.31 1.12 ;
        RECT  2.43 0.96 2.71 1.24 ;
        RECT  2.50 0.96 2.66 2.20 ;
        RECT  2.43 1.92 2.71 2.20 ;
        RECT  2.43 2.04 3.31 2.20 ;
        RECT  3.15 2.04 3.31 2.64 ;
        RECT  3.15 2.48 4.25 2.64 ;
        RECT  3.97 2.48 4.25 2.76 ;
        RECT  5.59 0.88 5.91 1.16 ;
        RECT  5.59 0.88 5.75 2.00 ;
        RECT  5.25 1.84 6.23 2.00 ;
        RECT  5.25 1.84 5.53 2.12 ;
        RECT  5.95 1.84 6.23 2.12 ;
        RECT  6.15 0.88 6.43 1.16 ;
        RECT  6.27 0.88 6.43 1.58 ;
        RECT  7.11 1.14 7.39 1.58 ;
        RECT  6.27 1.42 7.39 1.58 ;
        RECT  6.39 1.42 6.55 2.12 ;
        RECT  6.39 1.84 6.75 2.12 ;
        RECT  4.75 0.50 8.15 0.66 ;
        RECT  7.87 0.50 8.15 0.78 ;
        RECT  4.63 0.86 4.91 1.14 ;
        RECT  4.75 0.50 4.91 1.14 ;
        RECT  4.07 0.98 4.91 1.14 ;
        RECT  4.07 0.96 4.35 1.24 ;
        RECT  4.29 0.98 4.45 2.12 ;
        RECT  4.29 1.84 4.57 2.12 ;
        RECT  9.13 0.50 9.41 0.78 ;
        RECT  6.67 0.82 7.71 0.98 ;
        RECT  6.67 0.82 6.95 1.16 ;
        RECT  9.13 0.50 9.29 1.16 ;
        RECT  7.55 1.00 9.29 1.16 ;
        RECT  7.55 0.96 7.91 1.24 ;
        RECT  7.85 1.00 8.01 2.12 ;
        RECT  6.99 1.84 7.27 2.12 ;
        RECT  7.85 1.84 8.19 2.12 ;
        RECT  6.99 1.96 8.19 2.12 ;
        RECT  5.07 0.86 5.43 1.14 ;
        RECT  9.67 0.96 10.11 1.24 ;
        RECT  5.07 0.86 5.23 1.48 ;
        RECT  8.35 1.52 9.83 1.68 ;
        RECT  4.81 1.84 5.09 2.12 ;
        RECT  9.67 0.96 9.83 2.12 ;
        RECT  9.53 1.84 9.83 2.12 ;
        RECT  4.93 1.32 5.09 2.44 ;
        RECT  8.35 1.52 8.51 2.44 ;
        RECT  4.93 2.28 8.51 2.44 ;
        RECT  10.31 0.88 10.73 1.16 ;
        RECT  10.57 1.46 12.11 1.62 ;
        RECT  11.83 1.40 12.11 1.68 ;
        RECT  10.57 0.88 10.73 2.12 ;
        RECT  10.57 1.84 10.85 2.12 ;
        RECT  12.11 0.88 12.47 1.16 ;
        RECT  12.31 0.88 12.47 2.16 ;
        RECT  12.31 1.88 12.59 2.16 ;
        RECT  11.82 2.00 12.59 2.16 ;
        RECT  11.82 2.00 11.98 2.76 ;
        RECT  11.70 2.48 11.98 2.76 ;
    END
END DFFDERSSP8V1_0

MACRO DFFDERSSP4V1_0
    CLASS CORE ;
    FOREIGN DFFDERSSP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 30.02  LAYER ME1  ;
        ANTENNADIFFAREA 13.52  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.11  LAYER ME1  ;
        ANTENNAMAXAREACAR 26.95  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.55 1.46 13.94 1.74 ;
        RECT  13.43 1.90 13.71 2.50 ;
        RECT  13.55 0.64 13.71 2.50 ;
        RECT  13.43 0.64 13.71 1.24 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.66 0.44 11.94 0.94 ;
        RECT  11.45 0.44 11.94 0.72 ;
        END
    END SB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.99 1.40 10.41 1.68 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.24 1.40 3.54 1.76 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 29.65  LAYER ME1  ;
        ANTENNADIFFAREA 13.72  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.11  LAYER ME1  ;
        ANTENNAMAXAREACAR 26.63  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.88 1.19 2.32 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 2.04 1.19 2.32 ;
        RECT  0.91 0.88 1.19 1.16 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END E
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 30.02  LAYER ME1  ;
        ANTENNADIFFAREA 13.76  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.11  LAYER ME1  ;
        ANTENNAMAXAREACAR 26.95  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.47 1.90 14.75 2.50 ;
        RECT  14.47 0.64 14.75 1.24 ;
        RECT  14.47 0.64 14.74 2.50 ;
        RECT  14.46 1.46 14.74 1.74 ;
        END
    END QB
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 15.60 0.28 ;
        RECT  15.05 -0.28 15.42 0.32 ;
        RECT  14.99 0.64 15.27 1.24 ;
        RECT  15.05 -0.28 15.21 1.24 ;
        RECT  13.95 0.64 14.23 1.24 ;
        RECT  14.01 -0.28 14.17 1.24 ;
        RECT  12.91 0.64 13.19 1.24 ;
        RECT  12.97 -0.28 13.13 1.24 ;
        RECT  11.08 0.88 11.43 1.16 ;
        RECT  11.08 -0.28 11.24 1.16 ;
        RECT  8.69 -0.28 8.97 0.68 ;
        RECT  2.71 -0.28 2.99 0.64 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 15.60 3.48 ;
        RECT  15.05 2.88 15.42 3.48 ;
        RECT  14.99 1.90 15.27 2.50 ;
        RECT  15.05 1.90 15.21 3.48 ;
        RECT  13.95 1.90 14.23 2.50 ;
        RECT  14.01 1.90 14.17 3.48 ;
        RECT  12.91 1.90 13.19 2.50 ;
        RECT  12.97 1.90 13.13 3.48 ;
        RECT  12.31 2.40 12.59 3.48 ;
        RECT  11.09 1.84 11.37 2.12 ;
        RECT  11.15 1.84 11.31 3.48 ;
        RECT  10.05 1.84 10.33 2.12 ;
        RECT  10.11 1.84 10.27 3.48 ;
        RECT  8.77 1.96 9.29 2.12 ;
        RECT  9.01 1.84 9.29 2.12 ;
        RECT  8.65 2.52 8.93 3.48 ;
        RECT  8.77 1.96 8.93 3.48 ;
        RECT  2.71 2.52 2.99 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.95 0.88 2.23 1.16 ;
        RECT  1.95 2.04 2.23 2.32 ;
        RECT  2.07 0.88 2.23 2.70 ;
        RECT  2.07 2.42 2.37 2.70 ;
        RECT  2.27 0.44 2.55 0.72 ;
        RECT  1.55 0.56 2.55 0.72 ;
        RECT  1.55 0.56 1.71 1.16 ;
        RECT  1.43 0.88 1.71 1.16 ;
        RECT  1.49 0.88 1.65 2.32 ;
        RECT  1.43 2.04 1.71 2.32 ;
        RECT  3.47 0.96 3.86 1.24 ;
        RECT  3.70 1.46 4.02 1.74 ;
        RECT  3.70 0.96 3.86 2.20 ;
        RECT  3.47 1.92 3.86 2.20 ;
        RECT  4.07 0.44 4.35 0.72 ;
        RECT  3.15 0.56 4.35 0.72 ;
        RECT  3.15 0.56 3.31 1.12 ;
        RECT  2.43 0.96 3.31 1.12 ;
        RECT  2.43 0.96 2.71 1.24 ;
        RECT  2.50 0.96 2.66 2.20 ;
        RECT  2.43 1.92 2.71 2.20 ;
        RECT  2.43 2.04 3.31 2.20 ;
        RECT  3.15 2.04 3.31 2.64 ;
        RECT  3.15 2.48 4.25 2.64 ;
        RECT  3.97 2.48 4.25 2.76 ;
        RECT  5.59 0.88 5.91 1.16 ;
        RECT  5.59 0.88 5.75 2.00 ;
        RECT  5.25 1.84 6.23 2.00 ;
        RECT  5.25 1.84 5.53 2.12 ;
        RECT  5.95 1.84 6.23 2.12 ;
        RECT  6.15 0.88 6.43 1.16 ;
        RECT  6.27 0.88 6.43 1.58 ;
        RECT  7.11 1.14 7.39 1.58 ;
        RECT  6.27 1.42 7.39 1.58 ;
        RECT  6.39 1.42 6.55 2.12 ;
        RECT  6.39 1.84 6.75 2.12 ;
        RECT  4.75 0.50 8.15 0.66 ;
        RECT  7.87 0.50 8.15 0.78 ;
        RECT  4.63 0.86 4.91 1.14 ;
        RECT  4.75 0.50 4.91 1.14 ;
        RECT  4.07 0.98 4.91 1.14 ;
        RECT  4.07 0.96 4.35 1.24 ;
        RECT  4.29 0.98 4.45 2.12 ;
        RECT  4.29 1.84 4.57 2.12 ;
        RECT  9.13 0.50 9.41 0.78 ;
        RECT  6.67 0.82 7.71 0.98 ;
        RECT  6.67 0.82 6.95 1.16 ;
        RECT  9.13 0.50 9.29 1.16 ;
        RECT  7.55 1.00 9.29 1.16 ;
        RECT  7.55 0.96 7.91 1.24 ;
        RECT  7.85 1.00 8.01 2.12 ;
        RECT  6.99 1.84 7.27 2.12 ;
        RECT  7.85 1.84 8.19 2.12 ;
        RECT  6.99 1.96 8.19 2.12 ;
        RECT  5.07 0.86 5.43 1.14 ;
        RECT  9.67 0.96 10.11 1.24 ;
        RECT  5.07 0.86 5.23 1.48 ;
        RECT  8.35 1.52 9.83 1.68 ;
        RECT  4.81 1.84 5.09 2.12 ;
        RECT  9.67 0.96 9.83 2.12 ;
        RECT  9.53 1.84 9.83 2.12 ;
        RECT  4.93 1.32 5.09 2.44 ;
        RECT  8.35 1.52 8.51 2.44 ;
        RECT  4.93 2.28 8.51 2.44 ;
        RECT  10.31 0.88 10.73 1.16 ;
        RECT  10.57 1.46 12.11 1.62 ;
        RECT  11.83 1.40 12.11 1.68 ;
        RECT  10.57 0.88 10.73 2.12 ;
        RECT  10.57 1.84 10.85 2.12 ;
        RECT  12.11 0.88 12.47 1.16 ;
        RECT  12.31 0.88 12.47 2.16 ;
        RECT  12.31 1.88 12.59 2.16 ;
        RECT  11.82 2.00 12.59 2.16 ;
        RECT  11.82 2.00 11.98 2.76 ;
        RECT  11.70 2.48 11.98 2.76 ;
    END
END DFFDERSSP4V1_0

MACRO DFFDERSSP2V1_0
    CLASS CORE ;
    FOREIGN DFFDERSSP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 27.35  LAYER ME1  ;
        ANTENNADIFFAREA 12.38  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.83  LAYER ME1  ;
        ANTENNAMAXAREACAR 33.12  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.88 1.19 2.32 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 2.04 1.19 2.32 ;
        RECT  0.91 0.88 1.19 1.16 ;
        END
    END D
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 27.71  LAYER ME1  ;
        ANTENNADIFFAREA 12.17  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.83  LAYER ME1  ;
        ANTENNAMAXAREACAR 33.56  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.06 1.46 14.32 1.74 ;
        RECT  13.95 1.89 14.23 2.49 ;
        RECT  14.06 0.64 14.23 2.49 ;
        RECT  13.95 0.64 14.23 1.24 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 27.71  LAYER ME1  ;
        ANTENNADIFFAREA 12.17  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.83  LAYER ME1  ;
        ANTENNAMAXAREACAR 33.56  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.91 1.89 13.19 2.49 ;
        RECT  12.91 0.64 13.19 1.24 ;
        RECT  12.91 0.64 13.14 2.49 ;
        RECT  12.85 1.46 13.14 1.74 ;
        END
    END Q
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.99 1.40 10.41 1.68 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.24 1.40 3.54 1.76 ;
        END
    END CK
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.66 0.44 11.94 0.94 ;
        RECT  11.45 0.44 11.94 0.72 ;
        END
    END SB
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END E
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 14.40 3.48 ;
        RECT  13.94 2.88 14.22 3.48 ;
        RECT  13.43 1.89 13.71 2.49 ;
        RECT  13.49 1.89 13.65 3.48 ;
        RECT  12.31 2.40 12.59 3.48 ;
        RECT  11.09 1.84 11.37 2.12 ;
        RECT  11.15 1.84 11.31 3.48 ;
        RECT  10.05 1.84 10.33 2.12 ;
        RECT  10.11 1.84 10.27 3.48 ;
        RECT  8.77 1.96 9.29 2.12 ;
        RECT  9.01 1.84 9.29 2.12 ;
        RECT  8.65 2.52 8.93 3.48 ;
        RECT  8.77 1.96 8.93 3.48 ;
        RECT  2.71 2.52 2.99 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 14.40 0.28 ;
        RECT  13.94 -0.28 14.22 0.32 ;
        RECT  13.43 0.64 13.71 1.24 ;
        RECT  13.49 -0.28 13.65 1.24 ;
        RECT  11.08 0.88 11.43 1.16 ;
        RECT  11.08 -0.28 11.24 1.16 ;
        RECT  8.69 -0.28 8.97 0.68 ;
        RECT  2.71 -0.28 2.99 0.64 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.95 0.88 2.23 1.16 ;
        RECT  1.95 2.04 2.23 2.32 ;
        RECT  2.07 0.88 2.23 2.70 ;
        RECT  2.07 2.42 2.37 2.70 ;
        RECT  2.27 0.44 2.55 0.72 ;
        RECT  1.55 0.56 2.55 0.72 ;
        RECT  1.55 0.56 1.71 1.16 ;
        RECT  1.43 0.88 1.71 1.16 ;
        RECT  1.49 0.88 1.65 2.32 ;
        RECT  1.43 2.04 1.71 2.32 ;
        RECT  3.47 0.96 3.86 1.24 ;
        RECT  3.70 1.46 4.02 1.74 ;
        RECT  3.70 0.96 3.86 2.20 ;
        RECT  3.47 1.92 3.86 2.20 ;
        RECT  4.07 0.44 4.35 0.72 ;
        RECT  3.15 0.56 4.35 0.72 ;
        RECT  3.15 0.56 3.31 1.12 ;
        RECT  2.43 0.96 3.31 1.12 ;
        RECT  2.43 0.96 2.71 1.24 ;
        RECT  2.50 0.96 2.66 2.20 ;
        RECT  2.43 1.92 2.71 2.20 ;
        RECT  2.43 2.04 3.31 2.20 ;
        RECT  3.15 2.04 3.31 2.64 ;
        RECT  3.15 2.48 4.25 2.64 ;
        RECT  3.97 2.48 4.25 2.76 ;
        RECT  5.59 0.88 5.91 1.16 ;
        RECT  5.59 0.88 5.75 2.00 ;
        RECT  5.25 1.84 6.23 2.00 ;
        RECT  5.25 1.84 5.53 2.12 ;
        RECT  5.95 1.84 6.23 2.12 ;
        RECT  6.15 0.88 6.43 1.16 ;
        RECT  6.27 0.88 6.43 1.58 ;
        RECT  7.11 1.14 7.39 1.58 ;
        RECT  6.27 1.42 7.39 1.58 ;
        RECT  6.39 1.42 6.55 2.12 ;
        RECT  6.39 1.84 6.75 2.12 ;
        RECT  4.75 0.50 8.15 0.66 ;
        RECT  7.87 0.50 8.15 0.78 ;
        RECT  4.63 0.86 4.91 1.14 ;
        RECT  4.75 0.50 4.91 1.14 ;
        RECT  4.07 0.98 4.91 1.14 ;
        RECT  4.07 0.96 4.35 1.24 ;
        RECT  4.29 0.98 4.45 2.12 ;
        RECT  4.29 1.84 4.57 2.12 ;
        RECT  9.13 0.50 9.41 0.78 ;
        RECT  6.67 0.82 7.71 0.98 ;
        RECT  6.67 0.82 6.95 1.16 ;
        RECT  9.13 0.50 9.29 1.16 ;
        RECT  7.55 1.00 9.29 1.16 ;
        RECT  7.55 0.96 7.91 1.24 ;
        RECT  7.85 1.00 8.01 2.12 ;
        RECT  6.99 1.84 7.27 2.12 ;
        RECT  7.85 1.84 8.19 2.12 ;
        RECT  6.99 1.96 8.19 2.12 ;
        RECT  5.07 0.86 5.43 1.14 ;
        RECT  9.67 0.96 10.11 1.24 ;
        RECT  5.07 0.86 5.23 1.48 ;
        RECT  8.35 1.52 9.83 1.68 ;
        RECT  4.81 1.84 5.09 2.12 ;
        RECT  9.67 0.96 9.83 2.12 ;
        RECT  9.53 1.84 9.83 2.12 ;
        RECT  4.93 1.32 5.09 2.44 ;
        RECT  8.35 1.52 8.51 2.44 ;
        RECT  4.93 2.28 8.51 2.44 ;
        RECT  10.31 0.88 10.73 1.16 ;
        RECT  10.57 1.46 12.11 1.62 ;
        RECT  11.83 1.40 12.11 1.68 ;
        RECT  10.57 0.88 10.73 2.12 ;
        RECT  10.57 1.84 10.85 2.12 ;
        RECT  12.11 0.88 12.47 1.16 ;
        RECT  12.31 0.88 12.47 2.16 ;
        RECT  12.31 1.88 12.59 2.16 ;
        RECT  11.82 2.00 12.59 2.16 ;
        RECT  11.82 2.00 11.98 2.76 ;
        RECT  11.70 2.48 11.98 2.76 ;
    END
END DFFDERSSP2V1_0

MACRO DFFDERSSP1V1_0
    CLASS CORE ;
    FOREIGN DFFDERSSP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 27.26  LAYER ME1  ;
        ANTENNADIFFAREA 11.61  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER ME1  ;
        ANTENNAMAXAREACAR 40.56  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.88 1.19 2.32 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 2.04 1.19 2.32 ;
        RECT  0.91 0.88 1.19 1.16 ;
        END
    END D
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.66 0.44 11.94 0.94 ;
        RECT  11.45 0.44 11.94 0.72 ;
        END
    END SB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.24 1.40 3.54 1.76 ;
        END
    END CK
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.99 1.40 10.41 1.68 ;
        END
    END RB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 26.95  LAYER ME1  ;
        ANTENNADIFFAREA 11.41  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER ME1  ;
        ANTENNAMAXAREACAR 40.10  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.85 1.46 13.14 1.74 ;
        RECT  12.73 1.89 13.01 2.17 ;
        RECT  12.85 0.88 13.01 2.17 ;
        RECT  12.73 0.88 13.01 1.16 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 27.26  LAYER ME1  ;
        ANTENNADIFFAREA 11.41  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER ME1  ;
        ANTENNAMAXAREACAR 40.56  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.77 1.89 14.05 2.17 ;
        RECT  13.77 0.88 14.05 1.16 ;
        RECT  13.77 0.88 13.94 2.17 ;
        RECT  13.66 1.46 13.94 1.74 ;
        END
    END QB
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END E
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 14.40 0.28 ;
        RECT  13.94 -0.28 14.22 0.32 ;
        RECT  13.25 0.88 13.53 1.16 ;
        RECT  13.31 -0.28 13.47 1.16 ;
        RECT  11.08 0.88 11.43 1.16 ;
        RECT  11.08 -0.28 11.24 1.16 ;
        RECT  8.69 -0.28 8.97 0.68 ;
        RECT  2.71 -0.28 2.99 0.64 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 14.40 3.48 ;
        RECT  13.94 2.88 14.22 3.48 ;
        RECT  13.25 1.89 13.53 2.17 ;
        RECT  13.31 1.89 13.47 3.48 ;
        RECT  11.93 2.52 12.21 3.48 ;
        RECT  11.09 1.84 11.37 2.12 ;
        RECT  11.15 1.84 11.31 3.48 ;
        RECT  10.05 1.84 10.33 2.12 ;
        RECT  10.11 1.84 10.27 3.48 ;
        RECT  8.77 1.96 9.29 2.12 ;
        RECT  9.01 1.84 9.29 2.12 ;
        RECT  8.65 2.52 8.93 3.48 ;
        RECT  8.77 1.96 8.93 3.48 ;
        RECT  2.71 2.52 2.99 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.95 0.88 2.23 1.16 ;
        RECT  1.95 2.04 2.23 2.32 ;
        RECT  2.07 0.88 2.23 2.70 ;
        RECT  2.07 2.42 2.37 2.70 ;
        RECT  2.27 0.44 2.55 0.72 ;
        RECT  1.55 0.56 2.55 0.72 ;
        RECT  1.55 0.56 1.71 1.16 ;
        RECT  1.43 0.88 1.71 1.16 ;
        RECT  1.49 0.88 1.65 2.32 ;
        RECT  1.43 2.04 1.71 2.32 ;
        RECT  3.47 0.96 3.86 1.24 ;
        RECT  3.70 1.46 4.02 1.74 ;
        RECT  3.70 0.96 3.86 2.20 ;
        RECT  3.47 1.92 3.86 2.20 ;
        RECT  4.07 0.44 4.35 0.72 ;
        RECT  3.15 0.56 4.35 0.72 ;
        RECT  3.15 0.56 3.31 1.12 ;
        RECT  2.43 0.96 3.31 1.12 ;
        RECT  2.43 0.96 2.71 1.24 ;
        RECT  2.50 0.96 2.66 2.20 ;
        RECT  2.43 1.92 2.71 2.20 ;
        RECT  2.43 2.04 3.31 2.20 ;
        RECT  3.15 2.04 3.31 2.64 ;
        RECT  3.15 2.48 4.25 2.64 ;
        RECT  3.97 2.48 4.25 2.76 ;
        RECT  5.59 0.88 5.91 1.16 ;
        RECT  5.59 0.88 5.75 2.00 ;
        RECT  5.25 1.84 6.23 2.00 ;
        RECT  5.25 1.84 5.53 2.12 ;
        RECT  5.95 1.84 6.23 2.12 ;
        RECT  6.15 0.88 6.43 1.16 ;
        RECT  6.27 0.88 6.43 1.58 ;
        RECT  7.11 1.14 7.39 1.58 ;
        RECT  6.27 1.42 7.39 1.58 ;
        RECT  6.39 1.42 6.55 2.12 ;
        RECT  6.39 1.84 6.75 2.12 ;
        RECT  4.75 0.50 8.15 0.66 ;
        RECT  7.87 0.50 8.15 0.78 ;
        RECT  4.63 0.86 4.91 1.14 ;
        RECT  4.75 0.50 4.91 1.14 ;
        RECT  4.07 0.98 4.91 1.14 ;
        RECT  4.07 0.96 4.35 1.24 ;
        RECT  4.29 0.98 4.45 2.12 ;
        RECT  4.29 1.84 4.57 2.12 ;
        RECT  9.13 0.50 9.41 0.78 ;
        RECT  6.67 0.82 7.71 0.98 ;
        RECT  6.67 0.82 6.95 1.16 ;
        RECT  9.13 0.50 9.29 1.16 ;
        RECT  7.55 1.00 9.29 1.16 ;
        RECT  7.55 0.96 7.91 1.24 ;
        RECT  7.85 1.00 8.01 2.12 ;
        RECT  6.99 1.84 7.27 2.12 ;
        RECT  7.85 1.84 8.19 2.12 ;
        RECT  6.99 1.96 8.19 2.12 ;
        RECT  5.07 0.86 5.43 1.14 ;
        RECT  9.67 0.96 10.11 1.24 ;
        RECT  5.07 0.86 5.23 1.48 ;
        RECT  8.35 1.52 9.83 1.68 ;
        RECT  4.81 1.84 5.09 2.12 ;
        RECT  9.67 0.96 9.83 2.12 ;
        RECT  9.53 1.84 9.83 2.12 ;
        RECT  4.93 1.32 5.09 2.44 ;
        RECT  8.35 1.52 8.51 2.44 ;
        RECT  4.93 2.28 8.51 2.44 ;
        RECT  10.31 0.88 10.73 1.16 ;
        RECT  10.57 1.46 12.11 1.62 ;
        RECT  11.83 1.40 12.11 1.68 ;
        RECT  10.57 0.88 10.73 2.12 ;
        RECT  10.57 1.84 10.85 2.12 ;
        RECT  12.11 0.88 12.43 1.16 ;
        RECT  12.27 0.88 12.43 2.16 ;
        RECT  11.93 2.00 12.53 2.16 ;
        RECT  11.93 2.00 12.21 2.28 ;
        RECT  12.37 2.00 12.53 2.64 ;
        RECT  12.37 2.48 12.91 2.64 ;
        RECT  12.63 2.48 12.91 2.76 ;
    END
END DFFDERSSP1V1_0

MACRO DFFDERSP8V1_0
    CLASS CORE ;
    FOREIGN DFFDERSP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 31.57  LAYER ME1  ;
        ANTENNADIFFAREA 15.44  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.69  LAYER ME1  ;
        ANTENNAMAXAREACAR 18.68  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.91 1.90 15.19 2.50 ;
        RECT  14.91 0.64 15.19 1.24 ;
        RECT  14.91 0.64 15.07 2.50 ;
        RECT  13.99 1.52 15.07 1.68 ;
        RECT  13.99 1.46 14.34 1.74 ;
        RECT  13.87 1.90 14.15 2.50 ;
        RECT  13.99 0.64 14.15 2.50 ;
        RECT  13.87 0.64 14.15 1.24 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 31.57  LAYER ME1  ;
        ANTENNADIFFAREA 15.18  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.69  LAYER ME1  ;
        ANTENNAMAXAREACAR 18.68  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.83 1.90 13.11 2.50 ;
        RECT  12.83 0.64 13.11 1.24 ;
        RECT  12.83 0.64 12.99 2.50 ;
        RECT  11.91 1.52 12.99 1.68 ;
        RECT  11.91 1.46 12.34 1.74 ;
        RECT  11.79 1.90 12.07 2.50 ;
        RECT  11.91 0.64 12.07 2.50 ;
        RECT  11.79 0.64 12.07 1.24 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 31.57  LAYER ME1  ;
        ANTENNADIFFAREA 14.72  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.69  LAYER ME1  ;
        ANTENNAMAXAREACAR 18.68  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.81 1.19 2.25 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  0.91 0.81 1.19 1.09 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.22 1.40 3.54 1.76 ;
        END
    END CK
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.22 1.40 9.60 1.68 ;
        END
    END RB
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 16.00 0.28 ;
        RECT  15.49 -0.28 15.82 0.32 ;
        RECT  15.43 0.64 15.71 1.24 ;
        RECT  15.49 -0.28 15.65 1.24 ;
        RECT  14.39 0.64 14.67 1.24 ;
        RECT  14.45 -0.28 14.61 1.24 ;
        RECT  13.35 0.64 13.63 1.24 ;
        RECT  13.41 -0.28 13.57 1.24 ;
        RECT  12.31 0.64 12.59 1.24 ;
        RECT  12.37 -0.28 12.53 1.24 ;
        RECT  11.27 0.64 11.55 1.24 ;
        RECT  11.33 -0.28 11.49 1.24 ;
        RECT  10.27 0.88 10.55 1.16 ;
        RECT  10.33 -0.28 10.49 1.16 ;
        RECT  7.29 -0.28 7.57 0.72 ;
        RECT  2.71 -0.28 2.99 0.64 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 16.00 3.48 ;
        RECT  15.49 2.88 15.82 3.48 ;
        RECT  15.43 1.90 15.71 2.50 ;
        RECT  15.49 1.90 15.65 3.48 ;
        RECT  14.39 1.90 14.67 2.50 ;
        RECT  14.45 1.90 14.61 3.48 ;
        RECT  13.35 1.90 13.63 2.50 ;
        RECT  13.41 1.90 13.57 3.48 ;
        RECT  12.31 1.90 12.59 2.50 ;
        RECT  12.37 1.90 12.53 3.48 ;
        RECT  11.27 1.90 11.55 2.50 ;
        RECT  11.33 1.90 11.49 3.48 ;
        RECT  10.27 1.84 10.55 2.12 ;
        RECT  10.33 1.84 10.49 3.48 ;
        RECT  9.23 1.84 9.51 2.12 ;
        RECT  9.29 1.84 9.45 3.48 ;
        RECT  8.39 1.84 8.55 3.48 ;
        RECT  8.19 1.84 8.55 2.12 ;
        RECT  2.71 2.52 2.99 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.99 0.88 2.27 1.16 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.88 2.23 2.69 ;
        RECT  2.07 2.41 2.37 2.69 ;
        RECT  1.55 0.49 2.55 0.65 ;
        RECT  2.27 0.44 2.55 0.72 ;
        RECT  1.55 0.49 1.71 1.09 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  3.47 0.96 3.86 1.24 ;
        RECT  3.70 1.46 4.02 1.74 ;
        RECT  3.70 0.96 3.86 2.20 ;
        RECT  3.47 1.92 3.86 2.20 ;
        RECT  4.07 0.44 4.35 0.72 ;
        RECT  3.15 0.56 4.35 0.72 ;
        RECT  3.15 0.56 3.31 1.12 ;
        RECT  2.47 0.96 3.31 1.12 ;
        RECT  2.47 0.96 2.75 1.24 ;
        RECT  2.47 0.96 2.63 2.20 ;
        RECT  2.43 1.92 2.71 2.20 ;
        RECT  2.43 2.04 3.31 2.20 ;
        RECT  3.15 2.04 3.31 2.64 ;
        RECT  3.15 2.48 4.35 2.64 ;
        RECT  4.07 2.48 4.35 2.76 ;
        RECT  5.67 0.88 5.95 1.16 ;
        RECT  5.67 0.88 5.83 2.12 ;
        RECT  5.45 1.84 5.83 2.12 ;
        RECT  6.15 1.84 6.43 2.12 ;
        RECT  5.45 1.96 6.43 2.12 ;
        RECT  6.85 0.44 7.13 0.72 ;
        RECT  6.31 0.56 7.13 0.72 ;
        RECT  6.19 0.88 6.47 1.16 ;
        RECT  6.31 0.56 6.47 1.68 ;
        RECT  6.31 1.52 6.75 1.68 ;
        RECT  6.59 1.52 6.75 2.12 ;
        RECT  6.59 1.84 6.95 2.12 ;
        RECT  4.63 0.87 4.91 1.15 ;
        RECT  4.07 0.99 4.91 1.15 ;
        RECT  4.07 0.96 4.35 1.24 ;
        RECT  4.19 0.96 4.35 2.12 ;
        RECT  4.19 1.84 4.47 2.12 ;
        RECT  4.19 1.96 4.77 2.12 ;
        RECT  4.61 1.96 4.77 2.76 ;
        RECT  7.95 2.42 8.23 2.76 ;
        RECT  4.61 2.60 8.23 2.76 ;
        RECT  8.15 0.50 8.43 0.78 ;
        RECT  6.71 0.88 6.99 1.20 ;
        RECT  7.33 0.92 7.61 1.20 ;
        RECT  8.15 0.50 8.31 1.20 ;
        RECT  6.71 1.04 8.31 1.20 ;
        RECT  7.11 1.04 7.27 2.12 ;
        RECT  7.11 1.84 7.47 2.12 ;
        RECT  5.13 0.87 5.43 1.15 ;
        RECT  8.81 0.92 9.09 1.20 ;
        RECT  7.63 1.52 8.97 1.68 ;
        RECT  8.81 0.92 8.97 2.12 ;
        RECT  5.01 1.84 5.29 2.12 ;
        RECT  8.71 1.84 8.99 2.12 ;
        RECT  5.13 0.87 5.29 2.44 ;
        RECT  7.63 1.52 7.79 2.44 ;
        RECT  5.13 2.28 7.79 2.44 ;
        RECT  9.37 0.88 9.65 1.16 ;
        RECT  9.37 1.00 9.92 1.16 ;
        RECT  9.76 1.46 10.75 1.62 ;
        RECT  10.47 1.40 10.75 1.68 ;
        RECT  9.76 1.00 9.92 2.12 ;
        RECT  9.75 1.84 10.03 2.12 ;
        RECT  10.79 0.88 11.07 1.16 ;
        RECT  10.79 1.84 11.07 2.12 ;
        RECT  10.91 0.88 11.07 2.76 ;
        RECT  10.82 2.48 11.10 2.76 ;
    END
END DFFDERSP8V1_0

MACRO DFFDERSP4V1_0
    CLASS CORE ;
    FOREIGN DFFDERSP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 27.34  LAYER ME1  ;
        ANTENNADIFFAREA 12.40  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.11  LAYER ME1  ;
        ANTENNAMAXAREACAR 24.55  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.86 1.46 13.14 1.74 ;
        RECT  12.83 1.90 13.11 2.50 ;
        RECT  12.86 0.64 13.11 2.50 ;
        RECT  12.83 0.64 13.11 1.24 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 27.34  LAYER ME1  ;
        ANTENNADIFFAREA 12.14  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.11  LAYER ME1  ;
        ANTENNAMAXAREACAR 24.55  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.79 1.90 12.07 2.50 ;
        RECT  11.79 0.64 12.07 1.24 ;
        RECT  11.79 0.64 11.95 2.50 ;
        RECT  11.66 1.46 11.95 1.74 ;
        END
    END Q
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.22 1.40 9.60 1.68 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.22 1.40 3.54 1.76 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 27.34  LAYER ME1  ;
        ANTENNADIFFAREA 12.16  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.11  LAYER ME1  ;
        ANTENNAMAXAREACAR 24.55  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.81 1.19 2.25 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  0.91 0.81 1.19 1.09 ;
        END
    END D
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 14.00 0.28 ;
        RECT  13.41 -0.28 13.82 0.32 ;
        RECT  13.35 0.64 13.63 1.24 ;
        RECT  13.41 -0.28 13.57 1.24 ;
        RECT  12.31 0.64 12.59 1.24 ;
        RECT  12.37 -0.28 12.53 1.24 ;
        RECT  11.27 0.64 11.55 1.24 ;
        RECT  11.33 -0.28 11.49 1.24 ;
        RECT  10.27 0.88 10.55 1.16 ;
        RECT  10.33 -0.28 10.49 1.16 ;
        RECT  7.29 -0.28 7.57 0.72 ;
        RECT  2.71 -0.28 2.99 0.64 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 14.00 3.48 ;
        RECT  13.41 2.88 13.82 3.48 ;
        RECT  13.35 1.90 13.63 2.50 ;
        RECT  13.41 1.90 13.57 3.48 ;
        RECT  12.31 1.90 12.59 2.50 ;
        RECT  12.37 1.90 12.53 3.48 ;
        RECT  11.27 1.90 11.55 2.50 ;
        RECT  11.33 1.90 11.49 3.48 ;
        RECT  10.27 1.84 10.55 2.12 ;
        RECT  10.33 1.84 10.49 3.48 ;
        RECT  9.23 1.84 9.51 2.12 ;
        RECT  9.29 1.84 9.45 3.48 ;
        RECT  8.39 1.84 8.55 3.48 ;
        RECT  8.19 1.84 8.55 2.12 ;
        RECT  2.71 2.52 2.99 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.99 0.88 2.27 1.16 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.88 2.23 2.69 ;
        RECT  2.07 2.41 2.37 2.69 ;
        RECT  1.55 0.49 2.55 0.65 ;
        RECT  2.27 0.44 2.55 0.72 ;
        RECT  1.55 0.49 1.71 1.09 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  3.47 0.96 3.86 1.24 ;
        RECT  3.70 1.46 4.02 1.74 ;
        RECT  3.70 0.96 3.86 2.20 ;
        RECT  3.47 1.92 3.86 2.20 ;
        RECT  4.07 0.44 4.35 0.72 ;
        RECT  3.15 0.56 4.35 0.72 ;
        RECT  3.15 0.56 3.31 1.12 ;
        RECT  2.47 0.96 3.31 1.12 ;
        RECT  2.47 0.96 2.75 1.24 ;
        RECT  2.47 0.96 2.63 2.20 ;
        RECT  2.43 1.92 2.71 2.20 ;
        RECT  2.43 2.04 3.31 2.20 ;
        RECT  3.15 2.04 3.31 2.64 ;
        RECT  3.15 2.48 4.35 2.64 ;
        RECT  4.07 2.48 4.35 2.76 ;
        RECT  5.67 0.88 5.95 1.16 ;
        RECT  5.67 0.88 5.83 2.12 ;
        RECT  5.45 1.84 5.83 2.12 ;
        RECT  6.15 1.84 6.43 2.12 ;
        RECT  5.45 1.96 6.43 2.12 ;
        RECT  6.85 0.44 7.13 0.72 ;
        RECT  6.31 0.56 7.13 0.72 ;
        RECT  6.19 0.88 6.47 1.16 ;
        RECT  6.31 0.56 6.47 1.68 ;
        RECT  6.31 1.52 6.75 1.68 ;
        RECT  6.59 1.52 6.75 2.12 ;
        RECT  6.59 1.84 6.95 2.12 ;
        RECT  4.63 0.87 4.91 1.15 ;
        RECT  4.07 0.99 4.91 1.15 ;
        RECT  4.07 0.96 4.35 1.24 ;
        RECT  4.19 0.96 4.35 2.12 ;
        RECT  4.19 1.84 4.47 2.12 ;
        RECT  4.19 1.96 4.77 2.12 ;
        RECT  4.61 1.96 4.77 2.76 ;
        RECT  7.95 2.42 8.23 2.76 ;
        RECT  4.61 2.60 8.23 2.76 ;
        RECT  8.15 0.50 8.43 0.78 ;
        RECT  6.71 0.88 6.99 1.20 ;
        RECT  7.33 0.92 7.61 1.20 ;
        RECT  8.15 0.50 8.31 1.20 ;
        RECT  6.71 1.04 8.31 1.20 ;
        RECT  7.11 1.04 7.27 2.12 ;
        RECT  7.11 1.84 7.47 2.12 ;
        RECT  5.13 0.87 5.43 1.15 ;
        RECT  8.81 0.92 9.09 1.20 ;
        RECT  7.63 1.52 8.97 1.68 ;
        RECT  8.81 0.92 8.97 2.12 ;
        RECT  5.01 1.84 5.29 2.12 ;
        RECT  8.71 1.84 8.99 2.12 ;
        RECT  5.13 0.87 5.29 2.44 ;
        RECT  7.63 1.52 7.79 2.44 ;
        RECT  5.13 2.28 7.79 2.44 ;
        RECT  9.37 0.88 9.65 1.16 ;
        RECT  9.37 1.00 9.92 1.16 ;
        RECT  9.76 1.46 10.75 1.62 ;
        RECT  10.47 1.40 10.75 1.68 ;
        RECT  9.76 1.00 9.92 2.12 ;
        RECT  9.75 1.84 10.03 2.12 ;
        RECT  10.79 0.88 11.07 1.16 ;
        RECT  10.79 1.84 11.07 2.12 ;
        RECT  10.91 0.88 11.07 2.76 ;
        RECT  10.82 2.48 11.10 2.76 ;
    END
END DFFDERSP4V1_0

MACRO DFFDERSP2V1_0
    CLASS CORE ;
    FOREIGN DFFDERSP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 25.09  LAYER ME1  ;
        ANTENNADIFFAREA 10.82  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.83  LAYER ME1  ;
        ANTENNAMAXAREACAR 30.38  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.81 1.19 2.25 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  0.91 0.81 1.19 1.09 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.23 1.40 3.55 1.76 ;
        END
    END CK
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.22 1.40 9.60 1.68 ;
        END
    END RB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 25.09  LAYER ME1  ;
        ANTENNADIFFAREA 10.82  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.83  LAYER ME1  ;
        ANTENNAMAXAREACAR 30.38  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.27 1.90 11.55 2.50 ;
        RECT  11.27 0.64 11.55 1.24 ;
        RECT  11.27 0.64 11.54 2.50 ;
        RECT  11.26 1.46 11.54 1.74 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 25.09  LAYER ME1  ;
        ANTENNADIFFAREA 10.82  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.83  LAYER ME1  ;
        ANTENNAMAXAREACAR 30.38  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.43 1.46 12.72 1.74 ;
        RECT  12.31 1.90 12.59 2.50 ;
        RECT  12.43 0.64 12.59 2.50 ;
        RECT  12.31 0.64 12.59 1.24 ;
        END
    END QB
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 12.80 3.48 ;
        RECT  12.34 2.88 12.62 3.48 ;
        RECT  11.79 1.90 12.07 2.50 ;
        RECT  11.85 1.90 12.01 3.48 ;
        RECT  10.27 1.84 10.55 2.12 ;
        RECT  10.33 1.84 10.49 3.48 ;
        RECT  9.23 1.84 9.51 2.12 ;
        RECT  9.29 1.84 9.45 3.48 ;
        RECT  8.39 1.84 8.55 3.48 ;
        RECT  8.19 1.84 8.55 2.12 ;
        RECT  2.71 2.52 2.99 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 12.80 0.28 ;
        RECT  12.34 -0.28 12.62 0.32 ;
        RECT  11.79 0.64 12.07 1.24 ;
        RECT  11.85 -0.28 12.01 1.24 ;
        RECT  10.27 0.88 10.55 1.16 ;
        RECT  10.33 -0.28 10.49 1.16 ;
        RECT  7.29 -0.28 7.57 0.72 ;
        RECT  2.71 -0.28 2.99 0.64 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.99 0.88 2.27 1.16 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.88 2.23 2.69 ;
        RECT  2.07 2.41 2.37 2.69 ;
        RECT  1.55 0.49 2.55 0.65 ;
        RECT  2.27 0.44 2.55 0.72 ;
        RECT  1.55 0.49 1.71 1.09 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  3.47 0.96 3.87 1.24 ;
        RECT  3.71 1.46 4.03 1.74 ;
        RECT  3.71 0.96 3.87 2.20 ;
        RECT  3.47 1.92 3.87 2.20 ;
        RECT  4.07 0.44 4.35 0.72 ;
        RECT  3.15 0.56 4.35 0.72 ;
        RECT  3.15 0.56 3.31 1.12 ;
        RECT  2.47 0.96 3.31 1.12 ;
        RECT  2.47 0.96 2.75 1.24 ;
        RECT  2.47 0.96 2.63 2.20 ;
        RECT  2.43 1.92 2.71 2.20 ;
        RECT  2.43 2.04 3.31 2.20 ;
        RECT  3.15 2.04 3.31 2.64 ;
        RECT  3.15 2.48 4.35 2.64 ;
        RECT  4.07 2.48 4.35 2.76 ;
        RECT  5.67 0.88 5.95 1.16 ;
        RECT  5.67 0.88 5.83 2.12 ;
        RECT  5.45 1.84 5.83 2.12 ;
        RECT  6.15 1.84 6.43 2.12 ;
        RECT  5.45 1.96 6.43 2.12 ;
        RECT  6.85 0.44 7.13 0.72 ;
        RECT  6.31 0.56 7.13 0.72 ;
        RECT  6.19 0.88 6.47 1.16 ;
        RECT  6.31 0.56 6.47 1.68 ;
        RECT  6.31 1.52 6.75 1.68 ;
        RECT  6.59 1.52 6.75 2.12 ;
        RECT  6.59 1.84 6.95 2.12 ;
        RECT  4.63 0.87 4.91 1.15 ;
        RECT  4.07 0.99 4.91 1.15 ;
        RECT  4.07 0.96 4.35 1.24 ;
        RECT  4.19 0.96 4.35 2.12 ;
        RECT  4.19 1.84 4.47 2.12 ;
        RECT  4.19 1.96 4.77 2.12 ;
        RECT  4.61 1.96 4.77 2.76 ;
        RECT  7.95 2.42 8.23 2.76 ;
        RECT  4.61 2.60 8.23 2.76 ;
        RECT  8.15 0.50 8.43 0.78 ;
        RECT  6.71 0.88 6.99 1.20 ;
        RECT  7.33 0.92 7.61 1.20 ;
        RECT  8.15 0.50 8.31 1.20 ;
        RECT  6.71 1.04 8.31 1.20 ;
        RECT  7.11 1.04 7.27 2.12 ;
        RECT  7.11 1.84 7.47 2.12 ;
        RECT  5.13 0.87 5.43 1.15 ;
        RECT  8.81 0.92 9.09 1.20 ;
        RECT  7.63 1.52 8.97 1.68 ;
        RECT  8.81 0.92 8.97 2.12 ;
        RECT  5.01 1.84 5.29 2.12 ;
        RECT  8.71 1.84 8.99 2.12 ;
        RECT  5.13 0.87 5.29 2.44 ;
        RECT  7.63 1.52 7.79 2.44 ;
        RECT  5.13 2.28 7.79 2.44 ;
        RECT  9.37 0.88 9.65 1.16 ;
        RECT  9.37 1.00 9.92 1.16 ;
        RECT  9.76 1.46 10.75 1.62 ;
        RECT  10.47 1.40 10.75 1.68 ;
        RECT  9.76 1.00 9.92 2.12 ;
        RECT  9.75 1.84 10.03 2.12 ;
        RECT  10.79 0.88 11.07 1.16 ;
        RECT  10.79 1.84 11.07 2.12 ;
        RECT  10.91 0.88 11.07 2.76 ;
        RECT  10.82 2.48 11.10 2.76 ;
    END
END DFFDERSP2V1_0

MACRO DFFDERSP1V1_0
    CLASS CORE ;
    FOREIGN DFFDERSP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 24.36  LAYER ME1  ;
        ANTENNADIFFAREA 10.13  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER ME1  ;
        ANTENNAMAXAREACAR 36.24  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.43 1.46 12.72 1.74 ;
        RECT  12.31 1.90 12.59 2.18 ;
        RECT  12.43 0.88 12.59 2.18 ;
        RECT  12.31 0.88 12.59 1.16 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 24.67  LAYER ME1  ;
        ANTENNADIFFAREA 10.13  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER ME1  ;
        ANTENNAMAXAREACAR 36.71  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.27 1.90 11.55 2.18 ;
        RECT  11.27 0.88 11.55 1.16 ;
        RECT  11.27 0.88 11.54 2.18 ;
        RECT  11.26 1.46 11.54 1.74 ;
        END
    END Q
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.22 1.40 9.60 1.68 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.22 1.40 3.54 1.76 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 24.67  LAYER ME1  ;
        ANTENNADIFFAREA 10.13  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER ME1  ;
        ANTENNAMAXAREACAR 36.71  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.03 0.81 1.19 2.25 ;
        RECT  0.86 2.25 1.14 2.54 ;
        RECT  0.91 1.97 1.19 2.25 ;
        RECT  0.91 0.81 1.19 1.09 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.42 0.38 1.78 ;
        END
    END E
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 12.80 0.28 ;
        RECT  12.34 -0.28 12.62 0.32 ;
        RECT  11.79 0.88 12.07 1.16 ;
        RECT  11.85 -0.28 12.01 1.16 ;
        RECT  10.27 0.88 10.55 1.16 ;
        RECT  10.33 -0.28 10.49 1.16 ;
        RECT  7.29 -0.28 7.57 0.72 ;
        RECT  2.71 -0.28 2.99 0.64 ;
        RECT  0.32 -0.28 0.60 0.58 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 12.80 3.48 ;
        RECT  12.34 2.88 12.62 3.48 ;
        RECT  11.79 1.90 12.07 2.18 ;
        RECT  11.85 1.90 12.01 3.48 ;
        RECT  10.27 1.84 10.55 2.12 ;
        RECT  10.33 1.84 10.49 3.48 ;
        RECT  9.23 1.84 9.51 2.12 ;
        RECT  9.29 1.84 9.45 3.48 ;
        RECT  8.39 1.84 8.55 3.48 ;
        RECT  8.19 1.84 8.55 2.12 ;
        RECT  2.71 2.52 2.99 3.48 ;
        RECT  0.32 2.62 0.60 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.32 0.82 0.70 1.10 ;
        RECT  0.54 1.47 0.86 1.75 ;
        RECT  0.54 0.82 0.70 2.38 ;
        RECT  0.32 2.10 0.70 2.38 ;
        RECT  1.99 0.88 2.27 1.16 ;
        RECT  1.95 1.97 2.23 2.25 ;
        RECT  2.07 0.88 2.23 2.69 ;
        RECT  2.07 2.41 2.37 2.69 ;
        RECT  1.55 0.49 2.55 0.65 ;
        RECT  2.27 0.44 2.55 0.72 ;
        RECT  1.55 0.49 1.71 1.09 ;
        RECT  1.43 0.81 1.71 1.09 ;
        RECT  1.49 0.81 1.65 2.25 ;
        RECT  1.43 1.97 1.71 2.25 ;
        RECT  3.47 0.96 3.86 1.24 ;
        RECT  3.70 1.46 4.02 1.74 ;
        RECT  3.70 0.96 3.86 2.20 ;
        RECT  3.47 1.92 3.86 2.20 ;
        RECT  4.07 0.44 4.35 0.72 ;
        RECT  3.15 0.56 4.35 0.72 ;
        RECT  3.15 0.56 3.31 1.12 ;
        RECT  2.47 0.96 3.31 1.12 ;
        RECT  2.47 0.96 2.75 1.24 ;
        RECT  2.47 0.96 2.63 2.20 ;
        RECT  2.43 1.92 2.71 2.20 ;
        RECT  2.43 2.04 3.31 2.20 ;
        RECT  3.15 2.04 3.31 2.64 ;
        RECT  3.15 2.48 4.35 2.64 ;
        RECT  4.07 2.48 4.35 2.76 ;
        RECT  5.67 0.88 5.95 1.16 ;
        RECT  5.67 0.88 5.83 2.12 ;
        RECT  5.45 1.84 5.83 2.12 ;
        RECT  6.15 1.84 6.43 2.12 ;
        RECT  5.45 1.96 6.43 2.12 ;
        RECT  6.85 0.44 7.13 0.72 ;
        RECT  6.31 0.56 7.13 0.72 ;
        RECT  6.19 0.88 6.47 1.16 ;
        RECT  6.31 0.56 6.47 1.68 ;
        RECT  6.31 1.52 6.75 1.68 ;
        RECT  6.59 1.52 6.75 2.12 ;
        RECT  6.59 1.84 6.95 2.12 ;
        RECT  4.63 0.87 4.91 1.15 ;
        RECT  4.07 0.99 4.91 1.15 ;
        RECT  4.07 0.96 4.35 1.24 ;
        RECT  4.19 0.96 4.35 2.12 ;
        RECT  4.19 1.84 4.47 2.12 ;
        RECT  4.19 1.96 4.77 2.12 ;
        RECT  4.61 1.96 4.77 2.76 ;
        RECT  7.95 2.42 8.23 2.76 ;
        RECT  4.61 2.60 8.23 2.76 ;
        RECT  8.15 0.50 8.43 0.78 ;
        RECT  6.71 0.88 6.99 1.20 ;
        RECT  7.33 0.92 7.61 1.20 ;
        RECT  8.15 0.50 8.31 1.20 ;
        RECT  6.71 1.04 8.31 1.20 ;
        RECT  7.11 1.04 7.27 2.12 ;
        RECT  7.11 1.84 7.47 2.12 ;
        RECT  5.13 0.87 5.43 1.15 ;
        RECT  8.81 0.92 9.09 1.20 ;
        RECT  7.63 1.52 8.97 1.68 ;
        RECT  8.81 0.92 8.97 2.12 ;
        RECT  5.01 1.84 5.29 2.12 ;
        RECT  8.71 1.84 8.99 2.12 ;
        RECT  5.13 0.87 5.29 2.44 ;
        RECT  7.63 1.52 7.79 2.44 ;
        RECT  5.13 2.28 7.79 2.44 ;
        RECT  9.37 0.88 9.65 1.16 ;
        RECT  9.37 1.00 9.92 1.16 ;
        RECT  9.76 1.46 10.75 1.62 ;
        RECT  10.47 1.40 10.75 1.68 ;
        RECT  9.76 1.00 9.92 2.12 ;
        RECT  9.75 1.84 10.03 2.12 ;
        RECT  10.79 0.88 11.07 1.16 ;
        RECT  10.79 1.84 11.07 2.12 ;
        RECT  10.91 0.88 11.07 2.76 ;
        RECT  10.82 2.48 11.10 2.76 ;
    END
END DFFDERSP1V1_0

MACRO BUFSP8V1_0
    CLASS CORE ;
    FOREIGN BUFSP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.12  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.26 2.28 0.54 2.72 ;
        RECT  0.08 2.28 0.54 2.52 ;
        END
    END IN
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 5.53  LAYER ME1  ;
        ANTENNADIFFAREA 4.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.56  LAYER ME1  ;
        ANTENNAMAXAREACAR 9.93  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.26 1.84 2.54 2.12 ;
        RECT  2.26 0.96 2.54 1.24 ;
        RECT  2.26 0.96 2.42 2.12 ;
        RECT  1.32 1.52 2.42 1.68 ;
        RECT  1.22 1.84 1.50 2.12 ;
        RECT  1.22 0.96 1.50 1.24 ;
        RECT  1.32 0.96 1.48 2.12 ;
        END
    END OUT
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 3.20 0.28 ;
        RECT  2.78 0.66 3.06 0.94 ;
        RECT  2.74 -0.28 3.02 0.32 ;
        RECT  2.84 -0.28 3.00 0.94 ;
        RECT  1.74 0.66 2.02 0.94 ;
        RECT  1.80 -0.28 1.96 0.94 ;
        RECT  0.70 0.66 0.98 0.94 ;
        RECT  0.76 -0.28 0.92 0.94 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 3.20 3.48 ;
        RECT  2.78 2.14 3.06 2.42 ;
        RECT  2.74 2.88 3.02 3.48 ;
        RECT  2.84 2.14 3.00 3.48 ;
        RECT  1.74 2.14 2.02 2.42 ;
        RECT  1.80 2.14 1.96 3.48 ;
        RECT  0.70 2.14 0.98 2.42 ;
        RECT  0.76 2.14 0.92 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.96 0.38 1.24 ;
        RECT  0.20 1.46 1.16 1.62 ;
        RECT  0.88 1.40 1.16 1.68 ;
        RECT  0.20 0.96 0.36 2.12 ;
        RECT  0.14 1.84 0.42 2.12 ;
    END
END BUFSP8V1_0

MACRO BUFSP6V1_0
    CLASS CORE ;
    FOREIGN BUFSP6V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 2.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 4.79  LAYER ME1  ;
        ANTENNADIFFAREA 3.47  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.43  LAYER ME1  ;
        ANTENNAMAXAREACAR 11.08  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.26 1.84 2.54 2.12 ;
        RECT  2.26 0.96 2.54 1.24 ;
        RECT  2.26 0.96 2.42 2.12 ;
        RECT  1.32 1.52 2.42 1.68 ;
        RECT  1.22 1.84 1.50 2.12 ;
        RECT  1.22 0.96 1.50 1.24 ;
        RECT  1.32 0.96 1.48 2.12 ;
        END
    END OUT
    PIN IN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.12  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.26 2.28 0.54 2.72 ;
        RECT  0.08 2.28 0.54 2.52 ;
        END
    END IN
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 2.80 3.48 ;
        RECT  2.34 2.88 2.62 3.48 ;
        RECT  1.74 2.16 2.02 2.44 ;
        RECT  1.80 2.16 1.96 3.48 ;
        RECT  0.70 2.16 0.98 2.44 ;
        RECT  0.76 2.16 0.92 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 2.80 0.28 ;
        RECT  2.34 -0.28 2.62 0.32 ;
        RECT  1.74 0.64 2.02 0.92 ;
        RECT  1.80 -0.28 1.96 0.92 ;
        RECT  0.70 0.64 0.98 0.92 ;
        RECT  0.76 -0.28 0.92 0.92 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.96 0.38 1.24 ;
        RECT  0.20 1.46 1.16 1.62 ;
        RECT  0.88 1.40 1.16 1.68 ;
        RECT  0.20 0.96 0.36 2.12 ;
        RECT  0.14 1.84 0.42 2.12 ;
    END
END BUFSP6V1_0

MACRO BUFSP64V1_0
    CLASS CORE ;
    FOREIGN BUFSP64V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 27.61  LAYER ME1  ;
        ANTENNADIFFAREA 24.56  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 4.80  LAYER ME1  ;
        ANTENNAMAXAREACAR 5.75  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  15.28 1.84 15.56 2.12 ;
        RECT  15.28 0.96 15.56 1.24 ;
        RECT  15.28 0.96 15.44 2.12 ;
        RECT  2.92 1.52 15.44 1.68 ;
        RECT  14.24 1.84 14.52 2.12 ;
        RECT  14.24 0.96 14.52 1.24 ;
        RECT  14.30 0.96 14.46 2.12 ;
        RECT  13.20 1.84 13.48 2.12 ;
        RECT  13.20 0.96 13.48 1.24 ;
        RECT  13.26 0.96 13.42 2.12 ;
        RECT  12.14 1.84 12.42 2.12 ;
        RECT  12.14 0.96 12.42 1.24 ;
        RECT  12.20 0.96 12.36 2.12 ;
        RECT  11.10 1.84 11.38 2.12 ;
        RECT  11.10 0.96 11.38 1.24 ;
        RECT  11.16 0.96 11.32 2.12 ;
        RECT  10.06 1.84 10.34 2.12 ;
        RECT  10.06 0.96 10.34 1.24 ;
        RECT  10.12 0.96 10.28 2.12 ;
        RECT  9.02 1.84 9.30 2.12 ;
        RECT  9.02 0.96 9.30 1.24 ;
        RECT  9.08 0.96 9.24 2.12 ;
        RECT  7.98 1.84 8.26 2.12 ;
        RECT  7.98 0.96 8.26 1.24 ;
        RECT  8.04 0.96 8.20 2.12 ;
        RECT  6.94 1.84 7.22 2.12 ;
        RECT  6.94 0.96 7.22 1.24 ;
        RECT  7.00 0.96 7.16 2.12 ;
        RECT  5.90 1.84 6.18 2.12 ;
        RECT  5.90 0.96 6.18 1.24 ;
        RECT  5.96 0.96 6.12 2.12 ;
        RECT  4.86 1.84 5.14 2.12 ;
        RECT  4.86 0.96 5.14 1.24 ;
        RECT  4.92 0.96 5.08 2.12 ;
        RECT  3.82 1.84 4.10 2.12 ;
        RECT  3.82 0.96 4.10 1.24 ;
        RECT  3.88 0.96 4.04 2.12 ;
        RECT  2.78 1.84 3.08 2.12 ;
        RECT  2.92 0.96 3.08 2.12 ;
        RECT  2.78 0.96 3.08 1.24 ;
        END
    END OUT
    PIN IN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.71  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.40 0.60 1.68 ;
        RECT  0.08 1.40 0.34 1.74 ;
        END
    END IN
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 16.40 3.48 ;
        RECT  15.94 2.88 16.22 3.48 ;
        RECT  14.76 2.36 15.04 2.64 ;
        RECT  14.82 2.36 14.98 3.48 ;
        RECT  13.72 2.36 14.00 2.64 ;
        RECT  13.78 2.36 13.94 3.48 ;
        RECT  12.66 2.36 12.94 2.64 ;
        RECT  12.72 2.36 12.88 3.48 ;
        RECT  11.62 2.36 11.90 2.64 ;
        RECT  11.68 2.36 11.84 3.48 ;
        RECT  10.58 2.36 10.86 2.64 ;
        RECT  10.64 2.36 10.80 3.48 ;
        RECT  9.54 2.36 9.82 2.64 ;
        RECT  9.60 2.36 9.76 3.48 ;
        RECT  8.50 2.36 8.78 2.64 ;
        RECT  8.56 2.36 8.72 3.48 ;
        RECT  7.46 2.36 7.74 2.64 ;
        RECT  7.52 2.36 7.68 3.48 ;
        RECT  6.42 2.36 6.70 2.64 ;
        RECT  6.48 2.36 6.64 3.48 ;
        RECT  5.38 2.36 5.66 2.64 ;
        RECT  5.44 2.36 5.60 3.48 ;
        RECT  4.34 2.36 4.62 2.64 ;
        RECT  4.40 2.36 4.56 3.48 ;
        RECT  3.30 2.36 3.58 2.64 ;
        RECT  3.36 2.36 3.52 3.48 ;
        RECT  2.26 2.36 2.54 2.64 ;
        RECT  2.32 2.36 2.48 3.48 ;
        RECT  1.18 2.30 1.46 2.58 ;
        RECT  1.24 2.30 1.40 3.48 ;
        RECT  0.14 2.30 0.42 2.58 ;
        RECT  0.20 2.30 0.36 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 16.40 0.28 ;
        RECT  15.94 -0.28 16.22 0.32 ;
        RECT  14.76 0.44 15.04 0.72 ;
        RECT  14.82 -0.28 14.98 0.72 ;
        RECT  13.72 0.44 14.00 0.72 ;
        RECT  13.78 -0.28 13.94 0.72 ;
        RECT  12.66 0.44 12.94 0.72 ;
        RECT  12.72 -0.28 12.88 0.72 ;
        RECT  11.62 0.44 11.90 0.72 ;
        RECT  11.68 -0.28 11.84 0.72 ;
        RECT  10.58 0.44 10.86 0.72 ;
        RECT  10.64 -0.28 10.80 0.72 ;
        RECT  9.54 0.44 9.82 0.72 ;
        RECT  9.60 -0.28 9.76 0.72 ;
        RECT  8.50 0.44 8.78 0.72 ;
        RECT  8.56 -0.28 8.72 0.72 ;
        RECT  7.46 0.44 7.74 0.72 ;
        RECT  7.52 -0.28 7.68 0.72 ;
        RECT  6.42 0.44 6.70 0.72 ;
        RECT  6.48 -0.28 6.64 0.72 ;
        RECT  5.38 0.44 5.66 0.72 ;
        RECT  5.44 -0.28 5.60 0.72 ;
        RECT  4.34 0.44 4.62 0.72 ;
        RECT  4.40 -0.28 4.56 0.72 ;
        RECT  3.30 0.44 3.58 0.72 ;
        RECT  3.36 -0.28 3.52 0.72 ;
        RECT  2.26 0.44 2.54 0.72 ;
        RECT  2.32 -0.28 2.48 0.72 ;
        RECT  1.18 0.50 1.46 0.78 ;
        RECT  1.24 -0.28 1.40 0.78 ;
        RECT  0.14 0.50 0.42 0.78 ;
        RECT  0.20 -0.28 0.36 0.78 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.66 0.96 0.94 1.24 ;
        RECT  1.70 0.96 1.98 1.24 ;
        RECT  0.76 1.46 2.72 1.62 ;
        RECT  2.44 1.40 2.72 1.68 ;
        RECT  0.76 0.96 0.92 2.12 ;
        RECT  1.76 0.96 1.92 2.12 ;
        RECT  0.66 1.84 0.94 2.12 ;
        RECT  1.70 1.84 1.98 2.12 ;
    END
END BUFSP64V1_0

MACRO BUFSP4V1_0
    CLASS CORE ;
    FOREIGN BUFSP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 2.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 3.68  LAYER ME1  ;
        ANTENNADIFFAREA 2.54  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.31  LAYER ME1  ;
        ANTENNAMAXAREACAR 11.98  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.22 1.84 1.50 2.12 ;
        RECT  1.22 0.96 1.50 1.24 ;
        RECT  1.32 0.96 1.48 2.12 ;
        END
    END OUT
    PIN IN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 2.28 0.54 2.56 ;
        END
    END IN
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 2.40 3.48 ;
        RECT  1.80 2.88 2.22 3.48 ;
        RECT  1.74 2.20 2.02 2.48 ;
        RECT  1.80 2.20 1.96 3.48 ;
        RECT  0.70 2.20 0.98 2.48 ;
        RECT  0.76 2.20 0.92 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 2.40 0.28 ;
        RECT  1.80 -0.28 2.22 0.32 ;
        RECT  1.74 0.60 2.02 0.88 ;
        RECT  1.80 -0.28 1.96 0.88 ;
        RECT  0.70 0.60 0.98 0.88 ;
        RECT  0.76 -0.28 0.92 0.88 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.96 0.38 1.24 ;
        RECT  0.20 1.46 1.16 1.62 ;
        RECT  0.88 1.40 1.16 1.68 ;
        RECT  0.20 0.96 0.36 2.12 ;
        RECT  0.14 1.84 0.42 2.12 ;
    END
END BUFSP4V1_0

MACRO BUFSP48V1_0
    CLASS CORE ;
    FOREIGN BUFSP48V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.71  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.40 0.60 1.68 ;
        RECT  0.08 1.40 0.34 1.74 ;
        END
    END IN
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 21.49  LAYER ME1  ;
        ANTENNADIFFAREA 17.92  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 3.20  LAYER ME1  ;
        ANTENNAMAXAREACAR 6.72  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.06 1.84 11.34 2.12 ;
        RECT  11.06 0.96 11.34 1.24 ;
        RECT  11.06 0.96 11.22 2.12 ;
        RECT  2.86 1.52 11.22 1.68 ;
        RECT  10.02 1.84 10.30 2.12 ;
        RECT  10.02 0.96 10.30 1.24 ;
        RECT  10.08 0.96 10.24 2.12 ;
        RECT  8.98 1.84 9.26 2.12 ;
        RECT  8.98 0.96 9.26 1.24 ;
        RECT  9.04 0.96 9.20 2.12 ;
        RECT  7.94 1.84 8.22 2.12 ;
        RECT  7.94 0.96 8.22 1.24 ;
        RECT  8.00 0.96 8.16 2.12 ;
        RECT  6.90 1.84 7.18 2.12 ;
        RECT  6.90 0.96 7.18 1.24 ;
        RECT  6.96 0.96 7.12 2.12 ;
        RECT  5.86 1.84 6.14 2.12 ;
        RECT  5.86 0.96 6.14 1.24 ;
        RECT  5.92 0.96 6.08 2.12 ;
        RECT  4.82 1.84 5.10 2.12 ;
        RECT  4.82 0.96 5.10 1.24 ;
        RECT  4.88 0.96 5.04 2.12 ;
        RECT  3.78 1.84 4.06 2.12 ;
        RECT  3.78 0.96 4.06 1.24 ;
        RECT  3.84 0.96 4.00 2.12 ;
        RECT  2.74 1.84 3.02 2.12 ;
        RECT  2.86 0.96 3.02 2.12 ;
        RECT  2.74 0.96 3.02 1.24 ;
        END
    END OUT
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 12.80 0.28 ;
        RECT  12.34 -0.28 12.62 0.32 ;
        RECT  11.58 0.50 11.86 0.78 ;
        RECT  11.64 -0.28 11.80 0.78 ;
        RECT  10.54 0.50 10.82 0.78 ;
        RECT  10.60 -0.28 10.76 0.78 ;
        RECT  9.50 0.50 9.78 0.78 ;
        RECT  9.56 -0.28 9.72 0.78 ;
        RECT  8.46 0.50 8.74 0.78 ;
        RECT  8.52 -0.28 8.68 0.78 ;
        RECT  7.42 0.50 7.70 0.78 ;
        RECT  7.48 -0.28 7.64 0.78 ;
        RECT  6.38 0.50 6.66 0.78 ;
        RECT  6.44 -0.28 6.60 0.78 ;
        RECT  5.34 0.50 5.62 0.78 ;
        RECT  5.40 -0.28 5.56 0.78 ;
        RECT  4.30 0.50 4.58 0.78 ;
        RECT  4.36 -0.28 4.52 0.78 ;
        RECT  3.26 0.50 3.54 0.78 ;
        RECT  3.32 -0.28 3.48 0.78 ;
        RECT  2.22 0.50 2.50 0.78 ;
        RECT  2.28 -0.28 2.44 0.78 ;
        RECT  1.18 0.50 1.46 0.78 ;
        RECT  1.24 -0.28 1.40 0.78 ;
        RECT  0.14 0.50 0.42 0.78 ;
        RECT  0.20 -0.28 0.36 0.78 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 12.80 3.48 ;
        RECT  12.34 2.88 12.62 3.48 ;
        RECT  11.58 2.30 11.86 2.58 ;
        RECT  11.64 2.30 11.80 3.48 ;
        RECT  10.54 2.30 10.82 2.58 ;
        RECT  10.60 2.30 10.76 3.48 ;
        RECT  9.50 2.30 9.78 2.58 ;
        RECT  9.56 2.30 9.72 3.48 ;
        RECT  8.46 2.30 8.74 2.58 ;
        RECT  8.52 2.30 8.68 3.48 ;
        RECT  7.42 2.30 7.70 2.58 ;
        RECT  7.48 2.30 7.64 3.48 ;
        RECT  6.38 2.30 6.66 2.58 ;
        RECT  6.44 2.30 6.60 3.48 ;
        RECT  5.34 2.30 5.62 2.58 ;
        RECT  5.40 2.30 5.56 3.48 ;
        RECT  4.30 2.30 4.58 2.58 ;
        RECT  4.36 2.30 4.52 3.48 ;
        RECT  3.26 2.30 3.54 2.58 ;
        RECT  3.32 2.30 3.48 3.48 ;
        RECT  2.22 2.30 2.50 2.58 ;
        RECT  2.28 2.30 2.44 3.48 ;
        RECT  1.18 2.30 1.46 2.58 ;
        RECT  1.24 2.30 1.40 3.48 ;
        RECT  0.14 2.30 0.42 2.58 ;
        RECT  0.20 2.30 0.36 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.66 0.96 0.94 1.24 ;
        RECT  1.70 0.96 1.98 1.24 ;
        RECT  0.76 1.46 2.68 1.62 ;
        RECT  2.40 1.40 2.68 1.68 ;
        RECT  0.76 0.96 0.92 2.12 ;
        RECT  1.76 0.96 1.92 2.12 ;
        RECT  0.66 1.84 0.94 2.12 ;
        RECT  1.70 1.84 1.98 2.12 ;
    END
END BUFSP48V1_0

MACRO BUFSP3V1_0
    CLASS CORE ;
    FOREIGN BUFSP3V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 2.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 2.28 0.54 2.56 ;
        END
    END IN
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 3.78  LAYER ME1  ;
        ANTENNADIFFAREA 2.20  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.23  LAYER ME1  ;
        ANTENNAMAXAREACAR 16.42  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.22 1.84 1.50 2.12 ;
        RECT  1.22 0.96 1.50 1.24 ;
        RECT  1.32 0.96 1.48 2.12 ;
        END
    END OUT
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 2.40 0.28 ;
        RECT  1.80 -0.28 2.22 0.32 ;
        RECT  1.74 0.76 2.02 1.04 ;
        RECT  1.80 -0.28 1.96 1.04 ;
        RECT  0.70 0.76 0.98 1.04 ;
        RECT  0.76 -0.28 0.92 1.04 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 2.40 3.48 ;
        RECT  1.80 2.88 2.22 3.48 ;
        RECT  1.74 2.04 2.02 2.32 ;
        RECT  1.80 2.04 1.96 3.48 ;
        RECT  0.70 2.04 0.98 2.32 ;
        RECT  0.76 2.04 0.92 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.96 0.38 1.24 ;
        RECT  0.20 1.46 1.16 1.62 ;
        RECT  0.88 1.40 1.16 1.68 ;
        RECT  0.20 0.96 0.36 2.12 ;
        RECT  0.14 1.84 0.42 2.12 ;
    END
END BUFSP3V1_0

MACRO BUFSP32V1_0
    CLASS CORE ;
    FOREIGN BUFSP32V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.38  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.40 0.60 1.68 ;
        RECT  0.08 1.40 0.34 1.74 ;
        END
    END IN
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 13.94  LAYER ME1  ;
        ANTENNADIFFAREA 12.17  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.19  LAYER ME1  ;
        ANTENNAMAXAREACAR 6.37  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.94 1.84 7.22 2.12 ;
        RECT  6.94 0.96 7.22 1.24 ;
        RECT  6.94 0.96 7.10 2.12 ;
        RECT  1.84 1.52 7.10 1.68 ;
        RECT  5.90 1.84 6.18 2.12 ;
        RECT  5.90 0.96 6.18 1.24 ;
        RECT  5.96 0.96 6.12 2.12 ;
        RECT  4.86 1.84 5.14 2.12 ;
        RECT  4.86 0.96 5.14 1.24 ;
        RECT  4.92 0.96 5.08 2.12 ;
        RECT  3.82 1.84 4.10 2.12 ;
        RECT  3.82 0.96 4.10 1.24 ;
        RECT  3.88 0.96 4.04 2.12 ;
        RECT  2.78 1.84 3.06 2.12 ;
        RECT  2.78 0.96 3.06 1.24 ;
        RECT  2.84 0.96 3.00 2.12 ;
        RECT  1.74 1.84 2.02 2.12 ;
        RECT  1.74 0.96 2.02 1.24 ;
        RECT  1.84 0.96 2.00 2.12 ;
        END
    END OUT
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 8.40 0.28 ;
        RECT  7.94 -0.28 8.22 0.32 ;
        RECT  7.46 0.48 7.74 0.76 ;
        RECT  7.52 -0.28 7.68 0.76 ;
        RECT  6.42 0.48 6.70 0.76 ;
        RECT  6.48 -0.28 6.64 0.76 ;
        RECT  5.38 0.48 5.66 0.76 ;
        RECT  5.44 -0.28 5.60 0.76 ;
        RECT  4.34 0.48 4.62 0.76 ;
        RECT  4.40 -0.28 4.56 0.76 ;
        RECT  3.30 0.48 3.58 0.76 ;
        RECT  3.36 -0.28 3.52 0.76 ;
        RECT  2.26 0.48 2.54 0.76 ;
        RECT  2.32 -0.28 2.48 0.76 ;
        RECT  1.18 0.44 1.46 0.72 ;
        RECT  1.24 -0.28 1.40 0.72 ;
        RECT  0.14 0.44 0.42 0.72 ;
        RECT  0.20 -0.28 0.36 0.72 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 8.40 3.48 ;
        RECT  7.94 2.88 8.22 3.48 ;
        RECT  7.46 2.32 7.74 2.60 ;
        RECT  7.52 2.32 7.68 3.48 ;
        RECT  6.42 2.32 6.70 2.60 ;
        RECT  6.48 2.32 6.64 3.48 ;
        RECT  5.38 2.32 5.66 2.60 ;
        RECT  5.44 2.32 5.60 3.48 ;
        RECT  4.34 2.32 4.62 2.60 ;
        RECT  4.40 2.32 4.56 3.48 ;
        RECT  3.30 2.32 3.58 2.60 ;
        RECT  3.36 2.32 3.52 3.48 ;
        RECT  2.26 2.32 2.54 2.60 ;
        RECT  2.32 2.32 2.48 3.48 ;
        RECT  1.18 2.36 1.46 2.64 ;
        RECT  1.24 2.36 1.40 3.48 ;
        RECT  0.14 2.36 0.42 2.64 ;
        RECT  0.20 2.36 0.36 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.66 0.96 0.94 1.24 ;
        RECT  1.40 1.40 1.68 1.68 ;
        RECT  0.76 1.52 1.68 1.68 ;
        RECT  0.76 0.96 0.92 2.12 ;
        RECT  0.66 1.84 0.94 2.12 ;
    END
END BUFSP32V1_0

MACRO BUFSP2V1_0
    CLASS CORE ;
    FOREIGN BUFSP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 1.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.04  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 2.28 0.54 2.56 ;
        END
    END IN
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 2.52  LAYER ME1  ;
        ANTENNADIFFAREA 1.71  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.15  LAYER ME1  ;
        ANTENNAMAXAREACAR 16.94  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.22 1.84 1.50 2.12 ;
        RECT  1.22 0.96 1.50 1.24 ;
        RECT  1.32 0.96 1.48 2.12 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 1.60 3.48 ;
        RECT  1.14 2.88 1.42 3.48 ;
        RECT  0.70 2.18 0.98 2.46 ;
        RECT  0.76 2.18 0.92 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 1.60 0.28 ;
        RECT  1.14 -0.28 1.42 0.32 ;
        RECT  0.70 0.62 0.98 0.90 ;
        RECT  0.76 -0.28 0.92 0.90 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.90 0.38 1.18 ;
        RECT  0.22 1.46 1.16 1.62 ;
        RECT  0.88 1.40 1.16 1.68 ;
        RECT  0.22 0.90 0.38 2.12 ;
        RECT  0.10 1.84 0.38 2.12 ;
    END
END BUFSP2V1_0

MACRO BUFSP24V1_0
    CLASS CORE ;
    FOREIGN BUFSP24V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 11.72  LAYER ME1  ;
        ANTENNADIFFAREA 9.96  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.64  LAYER ME1  ;
        ANTENNAMAXAREACAR 7.14  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.90 1.84 6.18 2.12 ;
        RECT  5.90 0.96 6.18 1.24 ;
        RECT  5.90 0.96 6.06 2.12 ;
        RECT  1.84 1.52 6.06 1.68 ;
        RECT  4.86 1.84 5.14 2.12 ;
        RECT  4.86 0.96 5.14 1.24 ;
        RECT  4.92 0.96 5.08 2.12 ;
        RECT  3.82 1.84 4.10 2.12 ;
        RECT  3.82 0.96 4.10 1.24 ;
        RECT  3.88 0.96 4.04 2.12 ;
        RECT  2.78 1.84 3.06 2.12 ;
        RECT  2.78 0.96 3.06 1.24 ;
        RECT  2.84 0.96 3.00 2.12 ;
        RECT  1.74 1.84 2.02 2.12 ;
        RECT  1.74 0.96 2.02 1.24 ;
        RECT  1.84 0.96 2.00 2.12 ;
        END
    END OUT
    PIN IN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.38  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.32 1.40 0.60 1.68 ;
        RECT  0.08 1.48 0.48 1.72 ;
        END
    END IN
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 7.20 3.48 ;
        RECT  6.74 2.88 7.02 3.48 ;
        RECT  5.38 2.32 5.66 2.60 ;
        RECT  5.44 2.32 5.60 3.48 ;
        RECT  4.34 2.32 4.62 2.60 ;
        RECT  4.40 2.32 4.56 3.48 ;
        RECT  3.30 2.32 3.58 2.60 ;
        RECT  3.36 2.32 3.52 3.48 ;
        RECT  2.26 2.32 2.54 2.60 ;
        RECT  2.32 2.32 2.48 3.48 ;
        RECT  1.18 2.36 1.46 2.64 ;
        RECT  1.24 2.36 1.40 3.48 ;
        RECT  0.14 2.36 0.42 2.64 ;
        RECT  0.20 2.36 0.36 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 7.20 0.28 ;
        RECT  6.74 -0.28 7.02 0.32 ;
        RECT  5.38 0.48 5.66 0.76 ;
        RECT  5.44 -0.28 5.60 0.76 ;
        RECT  4.34 0.48 4.62 0.76 ;
        RECT  4.40 -0.28 4.56 0.76 ;
        RECT  3.30 0.48 3.58 0.76 ;
        RECT  3.36 -0.28 3.52 0.76 ;
        RECT  2.26 0.48 2.54 0.76 ;
        RECT  2.32 -0.28 2.48 0.76 ;
        RECT  1.18 0.44 1.46 0.72 ;
        RECT  1.24 -0.28 1.40 0.72 ;
        RECT  0.14 0.44 0.42 0.72 ;
        RECT  0.20 -0.28 0.36 0.72 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.66 0.96 0.94 1.24 ;
        RECT  1.40 1.40 1.68 1.68 ;
        RECT  0.76 1.52 1.68 1.68 ;
        RECT  0.76 0.96 0.92 2.12 ;
        RECT  0.66 1.84 0.94 2.12 ;
    END
END BUFSP24V1_0

MACRO BUFSP1V1_0
    CLASS CORE ;
    FOREIGN BUFSP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 1.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.40 0.74 1.74 ;
        END
    END IN
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 2.65  LAYER ME1  ;
        ANTENNADIFFAREA 1.25  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 39.48  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.14 1.90 1.48 2.18 ;
        RECT  1.32 0.58 1.48 2.18 ;
        RECT  1.14 0.58 1.48 0.86 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 1.60 3.48 ;
        RECT  1.14 2.88 1.42 3.48 ;
        RECT  0.62 1.90 0.90 2.18 ;
        RECT  0.68 1.90 0.84 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 1.60 0.28 ;
        RECT  1.14 -0.28 1.42 0.32 ;
        RECT  0.62 0.58 0.90 0.86 ;
        RECT  0.68 -0.28 0.84 0.86 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.08 0.58 0.38 0.86 ;
        RECT  0.08 1.08 1.16 1.24 ;
        RECT  0.88 1.04 1.16 1.32 ;
        RECT  0.08 0.58 0.24 2.18 ;
        RECT  0.08 1.90 0.38 2.18 ;
    END
END BUFSP1V1_0

MACRO BUFSP16V1_0
    CLASS CORE ;
    FOREIGN BUFSP16V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 9.14  LAYER ME1  ;
        ANTENNADIFFAREA 6.63  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.04  LAYER ME1  ;
        ANTENNAMAXAREACAR 8.78  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.82 1.84 5.10 2.12 ;
        RECT  4.82 0.96 5.10 1.24 ;
        RECT  4.82 0.96 4.98 2.12 ;
        RECT  1.80 1.52 4.98 1.68 ;
        RECT  3.78 1.84 4.06 2.12 ;
        RECT  3.78 0.96 4.06 1.24 ;
        RECT  3.84 0.96 4.00 2.12 ;
        RECT  2.74 1.84 3.02 2.12 ;
        RECT  2.74 0.96 3.02 1.24 ;
        RECT  2.80 0.96 2.96 2.12 ;
        RECT  1.70 1.84 1.98 2.12 ;
        RECT  1.70 0.96 1.98 1.24 ;
        RECT  1.80 0.96 1.96 2.12 ;
        END
    END OUT
    PIN IN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.23  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.40 0.56 1.68 ;
        RECT  0.08 1.40 0.34 1.74 ;
        END
    END IN
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 5.20 3.48 ;
        RECT  4.74 2.88 5.02 3.48 ;
        RECT  4.30 2.18 4.58 2.46 ;
        RECT  4.36 2.18 4.52 3.48 ;
        RECT  3.26 2.18 3.54 2.46 ;
        RECT  3.32 2.18 3.48 3.48 ;
        RECT  2.22 2.18 2.50 2.46 ;
        RECT  2.28 2.18 2.44 3.48 ;
        RECT  1.18 2.18 1.46 2.46 ;
        RECT  1.24 2.18 1.40 3.48 ;
        RECT  0.10 2.02 0.38 2.30 ;
        RECT  0.16 2.02 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 5.20 0.28 ;
        RECT  4.74 -0.28 5.02 0.32 ;
        RECT  4.30 0.62 4.58 0.90 ;
        RECT  4.36 -0.28 4.52 0.90 ;
        RECT  3.26 0.62 3.54 0.90 ;
        RECT  3.32 -0.28 3.48 0.90 ;
        RECT  2.22 0.62 2.50 0.90 ;
        RECT  2.28 -0.28 2.44 0.90 ;
        RECT  1.18 0.62 1.46 0.90 ;
        RECT  1.24 -0.28 1.40 0.90 ;
        RECT  0.10 0.74 0.38 1.02 ;
        RECT  0.16 -0.28 0.32 1.02 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.96 0.90 1.24 ;
        RECT  0.72 1.46 1.64 1.62 ;
        RECT  1.36 1.40 1.64 1.68 ;
        RECT  0.72 0.96 0.88 2.12 ;
        RECT  0.62 1.84 0.90 2.12 ;
    END
END BUFSP16V1_0

MACRO BUFSP12V1_0
    CLASS CORE ;
    FOREIGN BUFSP12V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.23  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.32 1.40 0.60 1.68 ;
        RECT  0.08 1.48 0.48 1.72 ;
        END
    END IN
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 7.54  LAYER ME1  ;
        ANTENNADIFFAREA 5.68  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.79  LAYER ME1  ;
        ANTENNAMAXAREACAR 9.52  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.88 1.84 4.16 2.12 ;
        RECT  3.88 0.96 4.16 1.24 ;
        RECT  3.88 0.96 4.04 2.12 ;
        RECT  1.84 1.52 4.04 1.68 ;
        RECT  2.78 1.84 3.06 2.12 ;
        RECT  2.78 0.96 3.06 1.24 ;
        RECT  2.84 0.96 3.00 2.12 ;
        RECT  1.74 1.84 2.02 2.12 ;
        RECT  1.74 0.96 2.02 1.24 ;
        RECT  1.84 0.96 2.00 2.12 ;
        END
    END OUT
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.40 0.28 ;
        RECT  3.94 -0.28 4.22 0.32 ;
        RECT  3.30 0.58 3.58 0.86 ;
        RECT  3.36 -0.28 3.52 0.86 ;
        RECT  2.26 0.58 2.54 0.86 ;
        RECT  2.32 -0.28 2.48 0.86 ;
        RECT  1.22 0.58 1.50 0.86 ;
        RECT  1.28 -0.28 1.44 0.86 ;
        RECT  0.10 0.74 0.38 1.02 ;
        RECT  0.16 -0.28 0.32 1.02 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.40 3.48 ;
        RECT  3.94 2.88 4.22 3.48 ;
        RECT  3.30 2.22 3.58 2.50 ;
        RECT  3.36 2.22 3.52 3.48 ;
        RECT  2.26 2.22 2.54 2.50 ;
        RECT  2.32 2.22 2.48 3.48 ;
        RECT  1.22 2.22 1.50 2.50 ;
        RECT  1.28 2.22 1.44 3.48 ;
        RECT  0.14 2.02 0.42 2.30 ;
        RECT  0.20 2.02 0.36 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.66 0.96 0.94 1.24 ;
        RECT  0.76 1.46 1.68 1.62 ;
        RECT  1.40 1.40 1.68 1.68 ;
        RECT  0.76 0.96 0.92 2.12 ;
        RECT  0.66 1.84 0.94 2.12 ;
    END
END BUFSP12V1_0

MACRO BUFCKSP8V1_0
    CLASS CORE ;
    FOREIGN BUFCKSP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.78  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.06 1.36 2.38 1.74 ;
        END
    END IN
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 10.77  LAYER ME1  ;
        ANTENNADIFFAREA 7.96  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.78  LAYER ME1  ;
        ANTENNAMAXAREACAR 13.85  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.74 1.98 6.10 2.14 ;
        RECT  5.82 1.86 6.10 2.14 ;
        RECT  4.82 0.92 5.10 1.20 ;
        RECT  4.78 1.86 5.06 2.14 ;
        RECT  4.82 0.92 4.98 2.14 ;
        RECT  3.90 1.46 4.34 1.74 ;
        RECT  3.74 1.86 4.06 2.14 ;
        RECT  3.90 0.92 4.06 2.14 ;
        RECT  3.78 0.92 4.06 1.20 ;
        END
    END OUT
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 7.20 0.28 ;
        RECT  6.74 -0.28 7.02 0.32 ;
        RECT  5.34 0.78 5.62 1.06 ;
        RECT  5.40 -0.28 5.56 1.06 ;
        RECT  4.30 0.78 4.58 1.06 ;
        RECT  4.36 -0.28 4.52 1.06 ;
        RECT  3.26 0.78 3.54 1.06 ;
        RECT  3.32 -0.28 3.48 1.06 ;
        RECT  2.22 0.78 2.50 1.06 ;
        RECT  2.28 -0.28 2.44 1.06 ;
        RECT  1.18 0.78 1.46 1.06 ;
        RECT  1.24 -0.28 1.40 1.06 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 7.20 3.48 ;
        RECT  6.74 2.88 7.02 3.48 ;
        RECT  6.34 2.38 6.62 2.66 ;
        RECT  6.40 2.38 6.56 3.48 ;
        RECT  5.30 2.38 5.58 2.66 ;
        RECT  5.36 2.38 5.52 3.48 ;
        RECT  4.26 2.38 4.54 2.66 ;
        RECT  4.32 2.38 4.48 3.48 ;
        RECT  3.22 2.38 3.50 2.66 ;
        RECT  3.28 2.38 3.44 3.48 ;
        RECT  2.18 2.38 2.46 2.66 ;
        RECT  2.24 2.38 2.40 3.48 ;
        RECT  1.14 2.38 1.42 2.66 ;
        RECT  1.20 2.38 1.36 3.48 ;
        RECT  0.10 2.38 0.38 2.66 ;
        RECT  0.16 2.38 0.32 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  1.70 0.92 1.98 1.20 ;
        RECT  2.74 0.92 3.02 1.20 ;
        RECT  3.42 1.40 3.72 1.68 ;
        RECT  1.70 0.92 1.86 2.14 ;
        RECT  0.62 1.86 1.94 2.02 ;
        RECT  2.70 1.86 3.58 2.02 ;
        RECT  3.42 1.40 3.58 2.02 ;
        RECT  0.62 1.86 0.90 2.14 ;
        RECT  2.82 0.92 2.98 2.14 ;
        RECT  1.66 1.98 2.98 2.14 ;
    END
END BUFCKSP8V1_0

MACRO BUFCKSP4V1_0
    CLASS CORE ;
    FOREIGN BUFCKSP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 6.02  LAYER ME1  ;
        ANTENNADIFFAREA 4.35  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.39  LAYER ME1  ;
        ANTENNAMAXAREACAR 15.49  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.18 1.98 3.50 2.14 ;
        RECT  3.22 1.86 3.50 2.14 ;
        RECT  2.34 1.46 2.74 1.74 ;
        RECT  2.18 1.86 2.50 2.14 ;
        RECT  2.34 0.92 2.50 2.14 ;
        RECT  2.22 0.92 2.50 1.20 ;
        END
    END OUT
    PIN IN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.39  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.82 1.36 1.14 1.74 ;
        END
    END IN
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.00 0.28 ;
        RECT  3.54 -0.28 3.82 0.32 ;
        RECT  2.74 0.78 3.02 1.06 ;
        RECT  2.80 -0.28 2.96 1.06 ;
        RECT  1.70 0.78 1.98 1.06 ;
        RECT  1.76 -0.28 1.92 1.06 ;
        RECT  0.66 0.78 0.94 1.06 ;
        RECT  0.72 -0.28 0.88 1.06 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.00 3.48 ;
        RECT  3.54 2.88 3.82 3.48 ;
        RECT  2.70 2.38 2.98 2.66 ;
        RECT  2.76 2.38 2.92 3.48 ;
        RECT  1.66 2.38 1.94 2.66 ;
        RECT  1.72 2.38 1.88 3.48 ;
        RECT  0.62 2.38 0.90 2.66 ;
        RECT  0.68 2.38 0.84 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  1.18 0.92 1.46 1.20 ;
        RECT  1.86 1.40 2.16 1.68 ;
        RECT  1.30 0.92 1.46 2.06 ;
        RECT  0.10 1.86 0.38 2.14 ;
        RECT  1.14 1.90 2.02 2.06 ;
        RECT  1.86 1.40 2.02 2.06 ;
        RECT  0.10 1.98 1.42 2.14 ;
        RECT  1.14 1.90 1.42 2.18 ;
    END
END BUFCKSP4V1_0

MACRO BUFCKSP3V1_0
    CLASS CORE ;
    FOREIGN BUFCKSP3V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.30  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.82 1.36 1.14 1.74 ;
        END
    END IN
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 5.29  LAYER ME1  ;
        ANTENNADIFFAREA 3.62  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.30  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.78  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.22 1.90 3.50 2.18 ;
        RECT  2.18 1.90 3.50 2.06 ;
        RECT  2.34 1.46 2.74 1.74 ;
        RECT  2.18 1.90 2.50 2.18 ;
        RECT  2.34 0.92 2.50 2.18 ;
        RECT  2.22 0.92 2.50 1.20 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 3.60 3.48 ;
        RECT  3.14 2.88 3.42 3.48 ;
        RECT  2.70 2.24 2.98 2.52 ;
        RECT  2.76 2.24 2.92 3.48 ;
        RECT  1.66 2.24 1.94 2.52 ;
        RECT  1.72 2.24 1.88 3.48 ;
        RECT  0.62 2.24 0.90 2.52 ;
        RECT  0.68 2.24 0.84 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 3.60 0.28 ;
        RECT  3.14 -0.28 3.42 0.32 ;
        RECT  1.70 0.58 1.98 0.86 ;
        RECT  1.76 -0.28 1.92 0.86 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  1.18 0.92 1.46 1.20 ;
        RECT  1.86 1.40 2.16 1.68 ;
        RECT  1.30 0.92 1.46 2.06 ;
        RECT  1.86 1.40 2.02 2.06 ;
        RECT  0.10 1.90 2.02 2.06 ;
        RECT  0.10 1.90 0.38 2.18 ;
        RECT  1.14 1.90 1.42 2.18 ;
    END
END BUFCKSP3V1_0

MACRO BUFCKSP32V1_0
    CLASS CORE ;
    FOREIGN BUFCKSP32V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 24.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 35.48  LAYER ME1  ;
        ANTENNADIFFAREA 27.88  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.96  LAYER ME1  ;
        ANTENNAMAXAREACAR 12.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.06 1.96 22.74 2.12 ;
        RECT  22.46 1.84 22.74 2.12 ;
        RECT  21.42 1.84 21.70 2.12 ;
        RECT  20.38 1.84 20.66 2.12 ;
        RECT  19.34 1.84 19.62 2.12 ;
        RECT  18.34 0.92 18.62 1.20 ;
        RECT  18.30 1.84 18.58 2.12 ;
        RECT  18.34 0.92 18.50 2.12 ;
        RECT  17.30 0.92 17.58 1.20 ;
        RECT  17.26 1.84 17.54 2.12 ;
        RECT  17.30 0.92 17.46 2.12 ;
        RECT  16.26 0.92 16.54 1.20 ;
        RECT  16.22 1.84 16.50 2.12 ;
        RECT  16.26 0.92 16.42 2.12 ;
        RECT  15.22 0.92 15.50 1.20 ;
        RECT  15.18 1.84 15.46 2.12 ;
        RECT  15.22 0.92 15.38 2.12 ;
        RECT  14.18 0.92 14.46 1.20 ;
        RECT  14.14 1.84 14.42 2.12 ;
        RECT  14.18 0.92 14.34 2.12 ;
        RECT  13.14 0.92 13.42 1.20 ;
        RECT  13.10 1.84 13.38 2.12 ;
        RECT  13.14 0.92 13.30 2.12 ;
        RECT  12.18 1.46 12.74 1.74 ;
        RECT  12.10 0.92 12.38 1.20 ;
        RECT  12.06 1.84 12.34 2.12 ;
        RECT  12.18 0.92 12.34 2.12 ;
        END
    END OUT
    PIN IN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.96  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.39 1.46 10.79 1.74 ;
        END
    END IN
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 24.00 0.28 ;
        RECT  23.54 -0.28 23.82 0.32 ;
        RECT  18.86 0.76 19.14 1.04 ;
        RECT  18.92 -0.28 19.08 1.04 ;
        RECT  17.82 0.76 18.10 1.04 ;
        RECT  17.88 -0.28 18.04 1.04 ;
        RECT  16.78 0.76 17.06 1.04 ;
        RECT  16.84 -0.28 17.00 1.04 ;
        RECT  15.74 0.76 16.02 1.04 ;
        RECT  15.80 -0.28 15.96 1.04 ;
        RECT  14.70 0.76 14.98 1.04 ;
        RECT  14.76 -0.28 14.92 1.04 ;
        RECT  13.66 0.76 13.94 1.04 ;
        RECT  13.72 -0.28 13.88 1.04 ;
        RECT  12.62 0.76 12.90 1.04 ;
        RECT  12.68 -0.28 12.84 1.04 ;
        RECT  11.58 0.76 11.86 1.04 ;
        RECT  11.64 -0.28 11.80 1.04 ;
        RECT  10.54 0.76 10.82 1.04 ;
        RECT  10.60 -0.28 10.76 1.04 ;
        RECT  9.50 0.76 9.78 1.04 ;
        RECT  9.56 -0.28 9.72 1.04 ;
        RECT  8.46 0.76 8.74 1.04 ;
        RECT  8.52 -0.28 8.68 1.04 ;
        RECT  7.42 0.76 7.70 1.04 ;
        RECT  7.48 -0.28 7.64 1.04 ;
        RECT  6.38 0.76 6.66 1.04 ;
        RECT  6.44 -0.28 6.60 1.04 ;
        RECT  5.34 0.76 5.62 1.04 ;
        RECT  5.40 -0.28 5.56 1.04 ;
        RECT  4.30 0.76 4.58 1.04 ;
        RECT  4.36 -0.28 4.52 1.04 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 24.00 3.48 ;
        RECT  23.54 2.88 23.82 3.48 ;
        RECT  22.98 2.40 23.26 2.68 ;
        RECT  23.04 2.40 23.20 3.48 ;
        RECT  21.94 2.40 22.22 2.68 ;
        RECT  22.00 2.40 22.16 3.48 ;
        RECT  20.90 2.40 21.18 2.68 ;
        RECT  20.96 2.40 21.12 3.48 ;
        RECT  19.86 2.40 20.14 2.68 ;
        RECT  19.92 2.40 20.08 3.48 ;
        RECT  18.82 2.40 19.10 2.68 ;
        RECT  18.88 2.40 19.04 3.48 ;
        RECT  17.78 2.40 18.06 2.68 ;
        RECT  17.84 2.40 18.00 3.48 ;
        RECT  16.74 2.40 17.02 2.68 ;
        RECT  16.80 2.40 16.96 3.48 ;
        RECT  15.70 2.40 15.98 2.68 ;
        RECT  15.76 2.40 15.92 3.48 ;
        RECT  14.66 2.40 14.94 2.68 ;
        RECT  14.72 2.40 14.88 3.48 ;
        RECT  13.62 2.40 13.90 2.68 ;
        RECT  13.68 2.40 13.84 3.48 ;
        RECT  12.58 2.40 12.86 2.68 ;
        RECT  12.64 2.40 12.80 3.48 ;
        RECT  11.54 2.40 11.82 2.68 ;
        RECT  11.60 2.40 11.76 3.48 ;
        RECT  10.50 2.40 10.78 2.68 ;
        RECT  10.56 2.40 10.72 3.48 ;
        RECT  9.46 2.40 9.74 2.68 ;
        RECT  9.52 2.40 9.68 3.48 ;
        RECT  8.42 2.40 8.70 2.68 ;
        RECT  8.48 2.40 8.64 3.48 ;
        RECT  7.38 2.40 7.66 2.68 ;
        RECT  7.44 2.40 7.60 3.48 ;
        RECT  6.34 2.40 6.62 2.68 ;
        RECT  6.40 2.40 6.56 3.48 ;
        RECT  5.30 2.40 5.58 2.68 ;
        RECT  5.36 2.40 5.52 3.48 ;
        RECT  4.26 2.40 4.54 2.68 ;
        RECT  4.32 2.40 4.48 3.48 ;
        RECT  3.22 2.40 3.50 2.68 ;
        RECT  3.28 2.40 3.44 3.48 ;
        RECT  2.18 2.40 2.46 2.68 ;
        RECT  2.24 2.40 2.40 3.48 ;
        RECT  1.14 2.40 1.42 2.68 ;
        RECT  1.20 2.40 1.36 3.48 ;
        RECT  0.10 2.40 0.38 2.68 ;
        RECT  0.16 2.40 0.32 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  4.82 0.92 5.10 1.20 ;
        RECT  5.86 0.92 6.14 1.20 ;
        RECT  6.90 0.92 7.18 1.20 ;
        RECT  7.94 0.92 8.22 1.20 ;
        RECT  8.98 0.92 9.26 1.20 ;
        RECT  10.02 0.92 10.30 1.20 ;
        RECT  11.06 0.92 11.34 1.20 ;
        RECT  11.74 1.40 12.02 1.68 ;
        RECT  4.82 0.92 4.98 2.12 ;
        RECT  5.86 0.92 6.02 2.12 ;
        RECT  6.90 0.92 7.06 2.12 ;
        RECT  7.94 0.92 8.10 2.12 ;
        RECT  8.98 0.92 9.14 2.12 ;
        RECT  10.02 0.92 10.18 2.12 ;
        RECT  11.02 1.89 11.90 2.05 ;
        RECT  0.62 1.84 10.26 2.00 ;
        RECT  11.74 1.40 11.90 2.05 ;
        RECT  0.62 1.84 0.90 2.12 ;
        RECT  1.66 1.84 1.94 2.12 ;
        RECT  2.70 1.84 2.98 2.12 ;
        RECT  3.74 1.84 4.02 2.12 ;
        RECT  4.78 1.84 5.06 2.12 ;
        RECT  5.82 1.84 6.10 2.12 ;
        RECT  6.86 1.84 7.14 2.12 ;
        RECT  7.90 1.84 8.18 2.12 ;
        RECT  8.94 1.84 9.22 2.12 ;
        RECT  9.98 1.96 11.30 2.12 ;
        RECT  11.14 0.92 11.30 2.17 ;
        RECT  11.02 1.89 11.30 2.17 ;
    END
END BUFCKSP32V1_0

MACRO BUFCKSP2V1_0
    CLASS CORE ;
    FOREIGN BUFCKSP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 2.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.16  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.36 1.18 1.74 ;
        END
    END IN
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 4.32  LAYER ME1  ;
        ANTENNADIFFAREA 2.35  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.16  LAYER ME1  ;
        ANTENNAMAXAREACAR 26.45  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.82 1.46 2.34 1.74 ;
        RECT  1.66 2.00 1.98 2.28 ;
        RECT  1.82 0.92 1.98 2.28 ;
        RECT  1.70 0.92 1.98 1.20 ;
        END
    END OUT
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 2.80 0.28 ;
        RECT  2.34 -0.28 2.62 0.32 ;
        RECT  1.18 0.88 1.46 1.16 ;
        RECT  1.24 -0.28 1.40 1.16 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 2.80 3.48 ;
        RECT  2.24 2.88 2.62 3.48 ;
        RECT  2.18 2.24 2.46 2.52 ;
        RECT  2.24 2.24 2.40 3.48 ;
        RECT  1.14 2.24 1.42 2.52 ;
        RECT  1.20 2.24 1.36 3.48 ;
        RECT  0.10 2.24 0.38 2.52 ;
        RECT  0.16 2.24 0.32 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.54 0.92 0.94 1.20 ;
        RECT  1.34 1.40 1.64 1.68 ;
        RECT  0.54 0.92 0.70 2.06 ;
        RECT  1.34 1.40 1.50 2.06 ;
        RECT  0.54 1.90 1.50 2.06 ;
        RECT  0.62 1.90 0.90 2.28 ;
    END
END BUFCKSP2V1_0

MACRO BUFCKSP1V1_0
    CLASS CORE ;
    FOREIGN BUFCKSP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 1.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 2.55  LAYER ME1  ;
        ANTENNADIFFAREA 1.73  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.10  LAYER ME1  ;
        ANTENNAMAXAREACAR 25.95  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.22 1.90 1.50 2.18 ;
        RECT  1.22 0.96 1.50 1.24 ;
        RECT  1.32 0.96 1.48 2.18 ;
        END
    END OUT
    PIN IN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.10  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.40 1.40 0.72 1.74 ;
        END
    END IN
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 1.60 3.48 ;
        RECT  1.14 2.88 1.42 3.48 ;
        RECT  0.70 2.28 0.98 2.56 ;
        RECT  0.76 2.28 0.92 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 1.60 0.28 ;
        RECT  1.14 -0.28 1.42 0.32 ;
        RECT  0.66 0.48 0.94 0.76 ;
        RECT  0.72 -0.28 0.88 0.76 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.08 0.96 0.38 1.24 ;
        RECT  0.88 1.46 1.16 1.74 ;
        RECT  0.08 0.96 0.24 2.18 ;
        RECT  0.88 1.46 1.04 2.06 ;
        RECT  0.08 1.90 1.04 2.06 ;
        RECT  0.08 1.90 0.46 2.18 ;
    END
END BUFCKSP1V1_0

MACRO BUFCKSP16V1_0
    CLASS CORE ;
    FOREIGN BUFCKSP16V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 18.28  LAYER ME1  ;
        ANTENNADIFFAREA 14.43  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.50  LAYER ME1  ;
        ANTENNAMAXAREACAR 12.22  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.34 1.96 11.82 2.12 ;
        RECT  11.54 1.84 11.82 2.12 ;
        RECT  10.50 1.84 10.78 2.12 ;
        RECT  9.50 0.92 9.78 1.20 ;
        RECT  9.46 1.84 9.74 2.12 ;
        RECT  9.50 0.92 9.66 2.12 ;
        RECT  8.46 0.92 8.74 1.20 ;
        RECT  8.42 1.84 8.70 2.12 ;
        RECT  8.46 0.92 8.62 2.12 ;
        RECT  7.42 0.92 7.70 1.20 ;
        RECT  7.38 1.84 7.66 2.12 ;
        RECT  7.42 0.92 7.58 2.12 ;
        RECT  6.46 1.46 6.74 1.74 ;
        RECT  6.38 0.92 6.66 1.20 ;
        RECT  6.34 1.84 6.62 2.12 ;
        RECT  6.46 0.92 6.62 2.12 ;
        END
    END OUT
    PIN IN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.50  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.84 1.46 5.24 1.74 ;
        END
    END IN
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 12.40 3.48 ;
        RECT  11.94 2.88 12.22 3.48 ;
        RECT  11.02 2.40 11.30 2.68 ;
        RECT  11.08 2.40 11.24 3.48 ;
        RECT  9.98 2.40 10.26 2.68 ;
        RECT  10.04 2.40 10.20 3.48 ;
        RECT  8.94 2.40 9.22 2.68 ;
        RECT  9.00 2.40 9.16 3.48 ;
        RECT  7.90 2.40 8.18 2.68 ;
        RECT  7.96 2.40 8.12 3.48 ;
        RECT  6.86 2.40 7.14 2.68 ;
        RECT  6.92 2.40 7.08 3.48 ;
        RECT  5.82 2.40 6.10 2.68 ;
        RECT  5.88 2.40 6.04 3.48 ;
        RECT  4.78 2.40 5.06 2.68 ;
        RECT  4.84 2.40 5.00 3.48 ;
        RECT  3.74 2.40 4.02 2.68 ;
        RECT  3.80 2.40 3.96 3.48 ;
        RECT  2.70 2.40 2.98 2.68 ;
        RECT  2.76 2.40 2.92 3.48 ;
        RECT  1.66 2.40 1.94 2.68 ;
        RECT  1.72 2.40 1.88 3.48 ;
        RECT  0.62 2.40 0.90 2.68 ;
        RECT  0.68 2.40 0.84 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 12.40 0.28 ;
        RECT  11.94 -0.28 12.22 0.32 ;
        RECT  8.98 0.74 9.26 1.02 ;
        RECT  9.04 -0.28 9.20 1.02 ;
        RECT  7.94 0.74 8.22 1.02 ;
        RECT  8.00 -0.28 8.16 1.02 ;
        RECT  6.90 0.74 7.18 1.02 ;
        RECT  6.96 -0.28 7.12 1.02 ;
        RECT  5.86 0.74 6.14 1.02 ;
        RECT  5.92 -0.28 6.08 1.02 ;
        RECT  4.82 0.74 5.10 1.02 ;
        RECT  4.88 -0.28 5.04 1.02 ;
        RECT  3.78 0.74 4.06 1.02 ;
        RECT  3.84 -0.28 4.00 1.02 ;
        RECT  2.74 0.74 3.02 1.02 ;
        RECT  2.80 -0.28 2.96 1.02 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  2.22 0.92 2.50 1.20 ;
        RECT  3.26 0.92 3.54 1.20 ;
        RECT  4.30 0.92 4.58 1.20 ;
        RECT  5.34 0.92 5.62 1.20 ;
        RECT  6.02 1.40 6.30 1.68 ;
        RECT  2.22 0.92 2.38 2.12 ;
        RECT  3.26 0.92 3.42 2.12 ;
        RECT  4.30 0.92 4.46 2.12 ;
        RECT  5.30 1.89 6.18 2.05 ;
        RECT  0.10 1.84 4.54 2.00 ;
        RECT  6.02 1.40 6.18 2.05 ;
        RECT  0.10 1.84 0.38 2.12 ;
        RECT  1.14 1.84 1.42 2.12 ;
        RECT  2.18 1.84 2.46 2.12 ;
        RECT  3.22 1.84 3.50 2.12 ;
        RECT  4.26 1.96 5.58 2.12 ;
        RECT  5.42 0.92 5.58 2.17 ;
        RECT  5.30 1.89 5.58 2.17 ;
    END
END BUFCKSP16V1_0

MACRO ANTSPV1_0
    CLASS CORE ;
    FOREIGN ANTSPV1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 0.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN
        DIRECTION INPUT ;
        ANTENNADIFFAREA 0.36  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAGATEAREA 0.00  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 0.64 0.70 1.24 ;
        END
    END IN
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 0.80 0.28 ;
        RECT  0.34 -0.28 0.62 0.32 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 0.80 3.48 ;
        RECT  0.34 2.88 0.62 3.48 ;
        END
    END VDD!
END ANTSPV1_0

MACRO AND4SP8V1_0
    CLASS CORE ;
    FOREIGN AND4SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 8.03  LAYER ME1  ;
        ANTENNADIFFAREA 5.99  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.58  LAYER ME1  ;
        ANTENNAMAXAREACAR 13.93  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.78 2.02 4.06 2.62 ;
        RECT  3.78 0.54 3.94 2.62 ;
        RECT  2.94 1.52 3.94 1.68 ;
        RECT  3.62 0.54 3.94 1.14 ;
        RECT  2.74 2.34 3.10 2.62 ;
        RECT  2.94 0.98 3.10 2.62 ;
        RECT  2.58 0.98 3.10 1.14 ;
        RECT  2.58 0.54 2.86 1.14 ;
        END
    END OUT
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.17  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.00 1.39 2.32 1.81 ;
        END
    END IN4
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.17  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.39 1.69 1.81 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.17  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.42 1.14 1.84 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.17  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.80 0.28 ;
        RECT  4.20 -0.28 4.62 0.32 ;
        RECT  4.14 0.54 4.42 1.14 ;
        RECT  4.20 -0.28 4.36 1.14 ;
        RECT  3.10 0.54 3.38 0.82 ;
        RECT  3.16 -0.28 3.32 0.82 ;
        RECT  2.02 0.44 2.30 1.14 ;
        RECT  2.08 -0.28 2.24 1.14 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.80 3.48 ;
        RECT  4.34 2.88 4.62 3.48 ;
        RECT  4.30 2.02 4.58 2.62 ;
        RECT  4.36 2.02 4.52 3.48 ;
        RECT  3.26 2.02 3.54 2.62 ;
        RECT  3.32 2.02 3.48 3.48 ;
        RECT  2.18 2.36 2.46 2.76 ;
        RECT  2.24 2.36 2.40 3.48 ;
        RECT  1.14 2.36 1.42 2.76 ;
        RECT  1.20 2.36 1.36 3.48 ;
        RECT  0.10 2.06 0.38 2.76 ;
        RECT  0.16 2.06 0.32 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.36 0.44 0.70 1.14 ;
        RECT  2.48 1.64 2.76 1.92 ;
        RECT  0.54 0.44 0.70 2.76 ;
        RECT  2.48 1.64 2.64 2.20 ;
        RECT  0.54 2.04 2.64 2.20 ;
        RECT  1.72 2.04 1.88 2.76 ;
        RECT  0.54 2.04 0.90 2.76 ;
        RECT  1.66 2.36 1.94 2.76 ;
    END
END AND4SP8V1_0

MACRO AND4SP4V1_0
    CLASS CORE ;
    FOREIGN AND4SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.14  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.14  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.14  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.39 1.69 1.81 ;
        END
    END IN3
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.14  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.00 1.39 2.32 1.81 ;
        END
    END IN4
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 6.63  LAYER ME1  ;
        ANTENNADIFFAREA 4.41  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.29  LAYER ME1  ;
        ANTENNAMAXAREACAR 23.02  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.74 2.34 3.10 2.62 ;
        RECT  2.94 0.98 3.10 2.62 ;
        RECT  2.92 1.52 3.10 1.68 ;
        RECT  2.58 0.98 3.10 1.14 ;
        RECT  2.58 0.54 2.86 1.14 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.00 3.48 ;
        RECT  3.32 2.88 3.82 3.48 ;
        RECT  3.26 2.02 3.54 2.62 ;
        RECT  3.32 2.02 3.48 3.48 ;
        RECT  2.18 2.34 2.46 2.74 ;
        RECT  2.24 2.34 2.40 3.48 ;
        RECT  1.14 2.34 1.42 2.74 ;
        RECT  1.20 2.34 1.36 3.48 ;
        RECT  0.10 2.16 0.38 2.74 ;
        RECT  0.16 2.16 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.00 0.28 ;
        RECT  3.54 -0.28 3.82 0.32 ;
        RECT  3.10 0.54 3.38 0.82 ;
        RECT  3.16 -0.28 3.32 0.82 ;
        RECT  2.02 0.50 2.30 1.08 ;
        RECT  2.08 -0.28 2.24 1.08 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.36 0.50 0.70 1.08 ;
        RECT  2.48 1.64 2.76 1.92 ;
        RECT  0.54 0.50 0.70 2.74 ;
        RECT  2.48 1.64 2.64 2.18 ;
        RECT  0.54 2.02 2.64 2.18 ;
        RECT  1.72 2.02 1.88 2.74 ;
        RECT  0.54 2.02 0.90 2.74 ;
        RECT  1.66 2.34 1.94 2.74 ;
    END
END AND4SP4V1_0

MACRO AND4SP2V1_0
    CLASS CORE ;
    FOREIGN AND4SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 5.26  LAYER ME1  ;
        ANTENNADIFFAREA 3.31  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.14  LAYER ME1  ;
        ANTENNAMAXAREACAR 36.49  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.74 2.34 3.10 2.62 ;
        RECT  2.94 0.54 3.10 2.62 ;
        RECT  2.92 1.52 3.10 1.68 ;
        RECT  2.58 0.54 3.10 1.14 ;
        END
    END OUT
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.10  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.00 1.39 2.32 1.81 ;
        END
    END IN4
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.10  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.39 1.69 1.81 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.10  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.10  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 3.20 0.28 ;
        RECT  2.74 -0.28 3.02 0.32 ;
        RECT  2.06 0.54 2.34 1.14 ;
        RECT  2.12 -0.28 2.28 1.14 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 3.20 3.48 ;
        RECT  2.74 2.88 3.02 3.48 ;
        RECT  2.18 2.34 2.46 2.74 ;
        RECT  2.24 2.34 2.40 3.48 ;
        RECT  1.14 2.34 1.42 2.74 ;
        RECT  1.20 2.34 1.36 3.48 ;
        RECT  0.10 2.34 0.38 2.74 ;
        RECT  0.16 2.34 0.32 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.36 0.68 0.64 1.08 ;
        RECT  2.48 1.64 2.76 1.92 ;
        RECT  2.48 1.64 2.64 2.18 ;
        RECT  0.54 2.02 2.64 2.18 ;
        RECT  0.54 0.80 0.70 2.74 ;
        RECT  1.72 2.02 1.88 2.74 ;
        RECT  0.54 2.34 0.90 2.74 ;
        RECT  1.66 2.34 1.94 2.74 ;
    END
END AND4SP2V1_0

MACRO AND4SP1V1_0
    CLASS CORE ;
    FOREIGN AND4SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.39 1.69 1.81 ;
        END
    END IN3
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 5.02  LAYER ME1  ;
        ANTENNADIFFAREA 2.43  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 74.63  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.70 2.34 3.10 2.62 ;
        RECT  2.94 0.80 3.10 2.62 ;
        RECT  2.92 1.52 3.10 1.68 ;
        RECT  2.54 0.80 3.10 1.08 ;
        END
    END OUT
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.06 1.39 2.34 1.81 ;
        END
    END IN4
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 3.20 0.28 ;
        RECT  2.74 -0.28 3.02 0.32 ;
        RECT  2.02 0.80 2.30 1.08 ;
        RECT  2.06 -0.28 2.22 1.08 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 3.20 3.48 ;
        RECT  2.74 2.88 3.02 3.48 ;
        RECT  2.18 2.34 2.46 2.62 ;
        RECT  2.24 2.34 2.40 3.48 ;
        RECT  1.14 2.34 1.42 2.62 ;
        RECT  1.20 2.34 1.36 3.48 ;
        RECT  0.10 2.34 0.38 2.62 ;
        RECT  0.16 2.34 0.32 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.36 0.80 0.70 1.08 ;
        RECT  2.50 1.90 2.78 2.18 ;
        RECT  0.54 2.02 2.78 2.18 ;
        RECT  0.54 0.80 0.70 2.62 ;
        RECT  1.66 2.02 1.82 2.62 ;
        RECT  0.54 2.34 0.90 2.62 ;
        RECT  1.66 2.34 1.94 2.62 ;
    END
END AND4SP1V1_0

MACRO AND4I1SP8V1_0
    CLASS CORE ;
    FOREIGN AND4I1SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.17  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.42 1.39 0.74 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.17  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.66 1.40 1.94 1.82 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.17  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.10 1.39 2.43 1.81 ;
        END
    END IN3
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 11.02  LAYER ME1  ;
        ANTENNADIFFAREA 7.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.74  LAYER ME1  ;
        ANTENNAMAXAREACAR 14.81  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.52 2.00 4.80 2.60 ;
        RECT  4.52 0.54 4.68 2.60 ;
        RECT  3.68 1.52 4.68 1.68 ;
        RECT  4.36 0.54 4.68 1.14 ;
        RECT  3.48 2.32 3.84 2.60 ;
        RECT  3.68 0.98 3.84 2.60 ;
        RECT  3.32 0.98 3.84 1.14 ;
        RECT  3.32 0.54 3.60 1.14 ;
        END
    END OUT
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.17  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.73 1.39 3.08 1.81 ;
        END
    END IN4
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 5.60 0.28 ;
        RECT  4.94 -0.28 5.42 0.32 ;
        RECT  4.88 0.54 5.16 1.14 ;
        RECT  4.94 -0.28 5.10 1.14 ;
        RECT  3.84 0.54 4.12 0.82 ;
        RECT  3.90 -0.28 4.06 0.82 ;
        RECT  2.76 0.44 3.04 1.14 ;
        RECT  2.81 -0.28 2.97 1.14 ;
        RECT  0.62 0.44 0.90 1.14 ;
        RECT  0.68 -0.28 0.84 1.14 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 5.60 3.48 ;
        RECT  5.10 2.88 5.42 3.48 ;
        RECT  5.04 2.00 5.32 2.60 ;
        RECT  5.10 2.00 5.26 3.48 ;
        RECT  4.00 2.00 4.28 2.60 ;
        RECT  4.06 2.00 4.22 3.48 ;
        RECT  2.92 2.34 3.20 2.74 ;
        RECT  2.98 2.34 3.14 3.48 ;
        RECT  1.88 2.34 2.16 2.74 ;
        RECT  1.94 2.34 2.10 3.48 ;
        RECT  0.84 2.34 1.12 2.74 ;
        RECT  0.90 2.34 1.06 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.44 0.38 1.14 ;
        RECT  0.90 1.38 1.18 1.66 ;
        RECT  0.90 1.38 1.06 2.13 ;
        RECT  0.10 1.97 1.06 2.13 ;
        RECT  0.10 0.44 0.26 2.74 ;
        RECT  0.10 2.34 0.60 2.74 ;
        RECT  1.10 0.44 1.50 1.14 ;
        RECT  3.24 1.53 3.52 1.81 ;
        RECT  3.24 1.53 3.40 2.16 ;
        RECT  1.34 2.00 3.40 2.16 ;
        RECT  1.34 0.44 1.50 2.74 ;
        RECT  2.40 2.00 2.56 2.74 ;
        RECT  1.34 2.34 1.64 2.74 ;
        RECT  2.40 2.34 2.68 2.74 ;
    END
END AND4I1SP8V1_0

MACRO AND4I1SP4V1_0
    CLASS CORE ;
    FOREIGN AND4I1SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.14  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.73 1.39 3.08 1.81 ;
        END
    END IN4
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 8.00  LAYER ME1  ;
        ANTENNADIFFAREA 5.17  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.43  LAYER ME1  ;
        ANTENNAMAXAREACAR 18.74  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.68 1.52 3.88 1.68 ;
        RECT  3.48 2.32 3.84 2.60 ;
        RECT  3.68 0.98 3.84 2.60 ;
        RECT  3.32 0.98 3.84 1.14 ;
        RECT  3.32 0.54 3.60 1.14 ;
        END
    END OUT
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.14  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.10 1.39 2.43 1.81 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.14  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.66 1.39 1.94 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.14  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.42 1.39 0.74 1.81 ;
        END
    END IN1
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.40 3.48 ;
        RECT  4.00 2.00 4.28 2.60 ;
        RECT  3.94 2.88 4.22 3.48 ;
        RECT  4.06 2.00 4.22 3.48 ;
        RECT  2.92 2.34 3.20 2.74 ;
        RECT  2.98 2.34 3.14 3.48 ;
        RECT  1.88 2.34 2.16 2.74 ;
        RECT  1.94 2.34 2.10 3.48 ;
        RECT  0.84 2.34 1.12 2.74 ;
        RECT  0.90 2.34 1.06 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.40 0.28 ;
        RECT  3.90 -0.28 4.22 0.32 ;
        RECT  3.84 0.54 4.12 0.82 ;
        RECT  3.90 -0.28 4.06 0.82 ;
        RECT  2.76 0.50 3.04 1.08 ;
        RECT  2.81 -0.28 2.97 1.08 ;
        RECT  0.62 0.50 0.90 1.08 ;
        RECT  0.68 -0.28 0.84 1.08 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.50 0.38 1.08 ;
        RECT  0.90 1.50 1.18 1.78 ;
        RECT  0.90 1.50 1.06 2.13 ;
        RECT  0.10 1.97 1.06 2.13 ;
        RECT  0.10 0.50 0.26 2.74 ;
        RECT  0.10 2.34 0.60 2.74 ;
        RECT  1.10 0.50 1.50 1.08 ;
        RECT  3.24 1.53 3.52 1.81 ;
        RECT  3.24 1.53 3.40 2.16 ;
        RECT  1.34 2.00 3.40 2.16 ;
        RECT  1.34 0.50 1.50 2.74 ;
        RECT  2.40 2.00 2.56 2.74 ;
        RECT  1.34 2.34 1.64 2.74 ;
        RECT  2.40 2.34 2.68 2.74 ;
    END
END AND4I1SP4V1_0

MACRO AND4I1SP2V1_0
    CLASS CORE ;
    FOREIGN AND4I1SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.10  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.42 1.39 0.74 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.10  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.66 1.39 1.94 1.81 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.10  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.10 1.39 2.43 1.81 ;
        END
    END IN3
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 7.09  LAYER ME1  ;
        ANTENNADIFFAREA 3.99  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.24  LAYER ME1  ;
        ANTENNAMAXAREACAR 29.56  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.48 2.38 3.88 2.66 ;
        RECT  3.72 0.54 3.88 2.66 ;
        RECT  3.32 0.54 3.88 1.14 ;
        END
    END OUT
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.10  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.73 1.39 3.12 1.81 ;
        END
    END IN4
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.00 0.28 ;
        RECT  3.54 -0.28 3.82 0.32 ;
        RECT  2.80 0.54 3.08 1.14 ;
        RECT  2.87 -0.28 3.03 1.14 ;
        RECT  0.62 0.68 0.90 1.08 ;
        RECT  0.68 -0.28 0.84 1.08 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.00 3.48 ;
        RECT  3.54 2.88 3.82 3.48 ;
        RECT  2.92 2.34 3.20 2.74 ;
        RECT  2.98 2.34 3.14 3.48 ;
        RECT  1.88 2.34 2.16 2.74 ;
        RECT  1.94 2.34 2.10 3.48 ;
        RECT  0.84 2.34 1.12 2.74 ;
        RECT  0.90 2.34 1.06 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.68 0.38 1.08 ;
        RECT  0.90 1.68 1.18 2.13 ;
        RECT  0.10 1.97 1.18 2.13 ;
        RECT  0.10 0.68 0.26 2.74 ;
        RECT  0.10 2.34 0.60 2.74 ;
        RECT  1.10 0.68 1.50 1.08 ;
        RECT  3.28 1.53 3.56 1.81 ;
        RECT  3.28 1.53 3.44 2.18 ;
        RECT  1.34 2.02 3.44 2.18 ;
        RECT  1.34 0.68 1.50 2.74 ;
        RECT  2.40 2.02 2.56 2.74 ;
        RECT  1.34 2.34 1.64 2.74 ;
        RECT  2.40 2.34 2.68 2.74 ;
    END
END AND4I1SP2V1_0

MACRO AND4I1SP1V1_0
    CLASS CORE ;
    FOREIGN AND4I1SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.73 1.39 3.14 1.81 ;
        END
    END IN4
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 6.72  LAYER ME1  ;
        ANTENNADIFFAREA 2.99  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        ANTENNAMAXAREACAR 49.99  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.44 2.34 3.88 2.62 ;
        RECT  3.72 0.80 3.88 2.62 ;
        RECT  3.28 0.80 3.88 1.08 ;
        END
    END OUT
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.10 1.39 2.43 1.81 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.66 1.39 1.94 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.42 1.39 0.74 1.81 ;
        END
    END IN1
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.00 3.48 ;
        RECT  3.54 2.88 3.82 3.48 ;
        RECT  2.92 2.34 3.20 2.62 ;
        RECT  2.98 2.34 3.14 3.48 ;
        RECT  1.88 2.34 2.16 2.62 ;
        RECT  1.94 2.34 2.10 3.48 ;
        RECT  0.84 2.34 1.12 2.62 ;
        RECT  0.90 2.34 1.06 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.00 0.28 ;
        RECT  3.54 -0.28 3.82 0.32 ;
        RECT  2.76 0.80 3.04 1.08 ;
        RECT  2.80 -0.28 2.96 1.08 ;
        RECT  0.62 0.80 0.90 1.08 ;
        RECT  0.68 -0.28 0.84 1.08 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.80 0.38 1.08 ;
        RECT  0.90 1.68 1.18 2.13 ;
        RECT  0.10 1.97 1.18 2.13 ;
        RECT  0.10 0.80 0.26 2.62 ;
        RECT  0.10 2.34 0.60 2.62 ;
        RECT  1.10 0.80 1.50 1.08 ;
        RECT  3.28 1.90 3.56 2.18 ;
        RECT  1.34 2.02 3.56 2.18 ;
        RECT  1.34 0.80 1.50 2.62 ;
        RECT  2.40 2.02 2.56 2.62 ;
        RECT  1.34 2.34 1.64 2.62 ;
        RECT  2.40 2.34 2.68 2.62 ;
    END
END AND4I1SP1V1_0

MACRO AND3SP8V1_0
    CLASS CORE ;
    FOREIGN AND3SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 8.42  LAYER ME1  ;
        ANTENNADIFFAREA 5.64  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.58  LAYER ME1  ;
        ANTENNAMAXAREACAR 14.62  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.26 2.02 3.54 2.62 ;
        RECT  3.26 0.54 3.42 2.62 ;
        RECT  2.26 1.52 3.42 1.68 ;
        RECT  3.14 0.54 3.42 1.14 ;
        RECT  2.22 2.02 2.50 2.62 ;
        RECT  2.26 0.54 2.42 2.62 ;
        RECT  2.10 0.54 2.42 1.14 ;
        END
    END OUT
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.17  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.17  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.17  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.46 1.62 1.81 ;
        END
    END IN3
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.40 3.48 ;
        RECT  3.84 2.88 4.22 3.48 ;
        RECT  3.78 2.02 4.06 2.62 ;
        RECT  3.84 2.02 4.00 3.48 ;
        RECT  2.74 2.02 3.02 2.62 ;
        RECT  2.80 2.02 2.96 3.48 ;
        RECT  1.66 2.48 1.94 2.76 ;
        RECT  1.72 2.48 1.88 3.48 ;
        RECT  0.62 2.48 0.90 2.76 ;
        RECT  0.68 2.48 0.84 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.40 0.28 ;
        RECT  3.72 -0.28 4.22 0.32 ;
        RECT  3.66 0.54 3.94 1.14 ;
        RECT  3.72 -0.28 3.88 1.14 ;
        RECT  2.62 0.54 2.90 1.14 ;
        RECT  2.68 -0.28 2.84 1.14 ;
        RECT  1.54 0.44 1.82 1.14 ;
        RECT  1.60 -0.28 1.76 1.14 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.26 0.44 0.70 1.14 ;
        RECT  1.82 1.46 2.10 1.74 ;
        RECT  0.54 0.44 0.70 2.18 ;
        RECT  1.82 1.46 1.98 2.18 ;
        RECT  0.12 2.02 1.98 2.18 ;
        RECT  0.12 2.02 0.28 2.62 ;
        RECT  1.14 2.02 1.30 2.62 ;
        RECT  0.10 2.34 0.38 2.62 ;
        RECT  1.14 2.34 1.42 2.62 ;
    END
END AND3SP8V1_0

MACRO AND3SP4V1_0
    CLASS CORE ;
    FOREIGN AND3SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.14  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.46 1.62 1.81 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.14  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.14  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 5.47  LAYER ME1  ;
        ANTENNADIFFAREA 3.76  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.29  LAYER ME1  ;
        ANTENNAMAXAREACAR 18.98  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.26 1.52 2.68 1.68 ;
        RECT  2.22 2.02 2.50 2.62 ;
        RECT  2.26 0.54 2.42 2.62 ;
        RECT  2.10 0.54 2.42 1.14 ;
        END
    END OUT
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 3.20 0.28 ;
        RECT  2.68 -0.28 3.02 0.32 ;
        RECT  2.62 0.54 2.90 1.14 ;
        RECT  2.68 -0.28 2.84 1.14 ;
        RECT  1.58 0.54 1.86 1.14 ;
        RECT  1.64 -0.28 1.80 1.14 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 3.20 3.48 ;
        RECT  2.74 2.88 3.02 3.48 ;
        RECT  2.74 2.02 3.02 2.62 ;
        RECT  2.80 2.02 2.96 3.48 ;
        RECT  1.66 2.48 1.94 2.76 ;
        RECT  1.72 2.48 1.88 3.48 ;
        RECT  0.62 2.48 0.90 2.76 ;
        RECT  0.68 2.48 0.84 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.26 0.54 0.70 1.12 ;
        RECT  1.82 1.46 2.10 1.74 ;
        RECT  0.54 0.54 0.70 2.18 ;
        RECT  1.82 1.46 1.98 2.18 ;
        RECT  0.12 2.02 1.98 2.18 ;
        RECT  0.12 2.02 0.28 2.62 ;
        RECT  1.14 2.02 1.30 2.62 ;
        RECT  0.10 2.34 0.38 2.62 ;
        RECT  1.14 2.34 1.42 2.62 ;
    END
END AND3SP4V1_0

MACRO AND3SP2V1_0
    CLASS CORE ;
    FOREIGN AND3SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 2.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 4.58  LAYER ME1  ;
        ANTENNADIFFAREA 2.89  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.14  LAYER ME1  ;
        ANTENNAMAXAREACAR 31.80  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.22 2.06 2.68 2.34 ;
        RECT  2.52 0.64 2.68 2.34 ;
        RECT  2.10 0.64 2.68 1.24 ;
        END
    END OUT
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.10  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.10  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.10  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.46 1.62 1.81 ;
        END
    END IN3
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 2.80 3.48 ;
        RECT  2.34 2.88 2.62 3.48 ;
        RECT  1.66 2.38 1.94 2.66 ;
        RECT  1.72 2.38 1.88 3.48 ;
        RECT  0.62 2.38 0.90 2.66 ;
        RECT  0.68 2.38 0.84 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 2.80 0.28 ;
        RECT  2.34 -0.28 2.62 0.32 ;
        RECT  1.58 0.64 1.86 1.24 ;
        RECT  1.64 -0.28 1.80 1.24 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.26 0.68 0.70 1.08 ;
        RECT  1.82 1.46 2.10 1.74 ;
        RECT  0.54 0.68 0.70 2.18 ;
        RECT  1.82 1.46 1.98 2.18 ;
        RECT  0.12 2.02 1.98 2.18 ;
        RECT  0.12 2.02 0.28 2.62 ;
        RECT  1.14 2.02 1.30 2.62 ;
        RECT  0.10 2.34 0.38 2.62 ;
        RECT  1.14 2.34 1.42 2.62 ;
    END
END AND3SP2V1_0

MACRO AND3SP1V1_0
    CLASS CORE ;
    FOREIGN AND3SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 2.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 4.39  LAYER ME1  ;
        ANTENNADIFFAREA 2.00  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 65.35  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.18 2.34 2.46 2.62 ;
        RECT  2.28 0.80 2.44 2.62 ;
        RECT  2.12 1.52 2.44 1.68 ;
        RECT  2.02 0.80 2.44 1.08 ;
        END
    END OUT
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.40 1.46 1.94 1.74 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.92 1.32 1.20 1.74 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.44 1.32 0.72 1.74 ;
        END
    END IN1
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 2.80 3.48 ;
        RECT  2.34 2.88 2.62 3.48 ;
        RECT  1.66 2.34 1.94 2.62 ;
        RECT  1.72 2.34 1.88 3.48 ;
        RECT  0.62 2.34 0.90 2.62 ;
        RECT  0.68 2.34 0.84 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 2.80 0.28 ;
        RECT  2.34 -0.28 2.62 0.32 ;
        RECT  1.50 0.80 1.78 1.08 ;
        RECT  1.54 -0.28 1.70 1.08 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.12 0.80 0.50 1.08 ;
        RECT  1.84 1.90 2.12 2.18 ;
        RECT  0.12 2.02 2.12 2.18 ;
        RECT  0.12 0.80 0.28 2.62 ;
        RECT  1.14 2.02 1.30 2.62 ;
        RECT  0.10 2.34 0.38 2.62 ;
        RECT  1.14 2.34 1.42 2.62 ;
    END
END AND3SP1V1_0

MACRO AND3OR2SP8V1_0
    CLASS CORE ;
    FOREIGN AND3OR2SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 11.83  LAYER ME1  ;
        ANTENNADIFFAREA 6.79  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.81  LAYER ME1  ;
        ANTENNAMAXAREACAR 14.59  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.24 2.04 5.52 2.64 ;
        RECT  5.24 0.56 5.52 1.16 ;
        RECT  5.30 0.56 5.46 2.64 ;
        RECT  4.52 1.52 5.46 1.68 ;
        RECT  4.20 2.04 4.68 2.20 ;
        RECT  4.52 1.00 4.68 2.20 ;
        RECT  4.20 1.00 4.68 1.16 ;
        RECT  4.20 2.04 4.48 2.32 ;
        RECT  4.20 0.56 4.48 1.16 ;
        END
    END OUT
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.17  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.26 1.39 3.59 1.81 ;
        END
    END IN4
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.40 1.46 1.94 1.74 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.92 1.32 1.20 1.74 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.44 1.32 0.72 1.74 ;
        END
    END IN1
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 6.40 0.28 ;
        RECT  5.82 -0.28 6.22 0.32 ;
        RECT  5.76 0.56 6.04 1.16 ;
        RECT  5.82 -0.28 5.98 1.16 ;
        RECT  4.72 0.56 5.00 0.84 ;
        RECT  4.78 -0.28 4.94 0.84 ;
        RECT  3.64 0.44 3.92 1.14 ;
        RECT  3.70 -0.28 3.86 1.14 ;
        RECT  2.60 0.44 2.88 0.72 ;
        RECT  2.66 -0.28 2.82 0.72 ;
        RECT  1.50 0.80 1.78 1.08 ;
        RECT  1.54 -0.28 1.70 1.08 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 6.40 3.48 ;
        RECT  5.82 2.88 6.22 3.48 ;
        RECT  5.76 2.04 6.04 2.64 ;
        RECT  5.82 2.04 5.98 3.48 ;
        RECT  4.72 2.36 5.00 2.64 ;
        RECT  4.78 2.36 4.94 3.48 ;
        RECT  3.64 2.48 3.92 2.76 ;
        RECT  3.70 2.48 3.86 3.48 ;
        RECT  1.66 2.34 1.94 2.62 ;
        RECT  1.72 2.34 1.88 3.48 ;
        RECT  0.62 2.34 0.90 2.62 ;
        RECT  0.68 2.34 0.84 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.12 0.80 0.50 1.08 ;
        RECT  1.84 1.90 2.12 2.18 ;
        RECT  0.12 2.02 2.12 2.18 ;
        RECT  0.12 0.80 0.28 2.62 ;
        RECT  1.14 2.02 1.30 2.62 ;
        RECT  0.10 2.34 0.38 2.62 ;
        RECT  1.14 2.34 1.42 2.62 ;
        RECT  2.02 0.80 2.44 1.08 ;
        RECT  2.28 1.46 2.78 1.74 ;
        RECT  2.28 0.80 2.44 2.62 ;
        RECT  2.18 2.34 2.46 2.62 ;
        RECT  3.12 0.68 3.40 0.96 ;
        RECT  3.12 0.68 3.28 1.23 ;
        RECT  2.94 1.07 3.28 1.23 ;
        RECT  3.82 1.46 4.10 1.74 ;
        RECT  2.94 1.97 3.98 2.13 ;
        RECT  3.82 1.46 3.98 2.13 ;
        RECT  2.94 1.07 3.10 2.76 ;
        RECT  2.74 2.06 3.10 2.76 ;
    END
END AND3OR2SP8V1_0

MACRO AND3OR2SP4V1_0
    CLASS CORE ;
    FOREIGN AND3OR2SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.44 1.32 0.72 1.74 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.92 1.32 1.20 1.74 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.40 1.46 1.94 1.74 ;
        END
    END IN3
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.14  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.26 1.39 3.54 1.81 ;
        END
    END IN4
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 9.01  LAYER ME1  ;
        ANTENNADIFFAREA 5.03  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER ME1  ;
        ANTENNAMAXAREACAR 18.23  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.20 2.04 4.68 2.20 ;
        RECT  4.52 1.00 4.68 2.20 ;
        RECT  4.20 1.00 4.68 1.16 ;
        RECT  4.20 2.04 4.48 2.32 ;
        RECT  4.20 0.56 4.48 1.16 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 5.20 3.48 ;
        RECT  4.74 2.88 5.02 3.48 ;
        RECT  4.72 2.36 5.00 2.64 ;
        RECT  4.78 2.36 4.94 3.48 ;
        RECT  3.64 2.48 3.92 2.76 ;
        RECT  3.70 2.48 3.86 3.48 ;
        RECT  1.66 2.34 1.94 2.62 ;
        RECT  1.72 2.34 1.88 3.48 ;
        RECT  0.62 2.34 0.90 2.62 ;
        RECT  0.68 2.34 0.84 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 5.20 0.28 ;
        RECT  4.74 -0.28 5.02 0.32 ;
        RECT  4.72 0.56 5.00 0.84 ;
        RECT  4.78 -0.28 4.94 0.84 ;
        RECT  3.68 0.56 3.96 1.16 ;
        RECT  3.74 -0.28 3.90 1.16 ;
        RECT  2.60 0.56 2.88 0.84 ;
        RECT  2.66 -0.28 2.82 0.84 ;
        RECT  1.50 0.80 1.78 1.08 ;
        RECT  1.54 -0.28 1.70 1.08 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.12 0.80 0.50 1.08 ;
        RECT  1.84 1.90 2.12 2.18 ;
        RECT  0.12 2.02 2.12 2.18 ;
        RECT  0.12 0.80 0.28 2.62 ;
        RECT  1.14 2.02 1.30 2.62 ;
        RECT  0.10 2.34 0.38 2.62 ;
        RECT  1.14 2.34 1.42 2.62 ;
        RECT  2.02 0.80 2.44 1.08 ;
        RECT  2.28 1.46 2.78 1.74 ;
        RECT  2.28 0.80 2.44 2.62 ;
        RECT  2.18 2.34 2.46 2.62 ;
        RECT  3.12 0.68 3.40 0.96 ;
        RECT  3.12 0.68 3.28 1.23 ;
        RECT  2.94 1.07 3.28 1.23 ;
        RECT  3.82 1.46 4.10 1.74 ;
        RECT  3.82 1.46 3.98 2.13 ;
        RECT  2.94 1.97 3.98 2.13 ;
        RECT  2.94 1.07 3.10 2.76 ;
        RECT  2.74 2.18 3.10 2.76 ;
    END
END AND3OR2SP4V1_0

MACRO AND3OR2SP2V1_0
    CLASS CORE ;
    FOREIGN AND3OR2SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 8.29  LAYER ME1  ;
        ANTENNADIFFAREA 4.11  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.31  LAYER ME1  ;
        ANTENNAMAXAREACAR 26.99  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.20 2.06 4.68 2.22 ;
        RECT  4.52 0.98 4.68 2.22 ;
        RECT  4.20 0.98 4.68 1.14 ;
        RECT  4.20 2.06 4.48 2.34 ;
        RECT  4.20 0.54 4.48 1.14 ;
        END
    END OUT
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.10  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.26 1.39 3.54 1.81 ;
        END
    END IN4
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.40 1.46 1.94 1.74 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.92 1.32 1.20 1.74 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.44 1.32 0.72 1.74 ;
        END
    END IN1
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.80 0.28 ;
        RECT  4.34 -0.28 4.62 0.32 ;
        RECT  3.68 0.54 3.96 1.14 ;
        RECT  3.74 -0.28 3.90 1.14 ;
        RECT  2.60 0.54 2.88 0.82 ;
        RECT  2.66 -0.28 2.82 0.82 ;
        RECT  1.50 0.80 1.78 1.08 ;
        RECT  1.54 -0.28 1.70 1.08 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.80 3.48 ;
        RECT  4.34 2.88 4.62 3.48 ;
        RECT  3.68 2.38 3.96 2.66 ;
        RECT  3.74 2.38 3.90 3.48 ;
        RECT  1.66 2.34 1.94 2.62 ;
        RECT  1.72 2.34 1.88 3.48 ;
        RECT  0.62 2.34 0.90 2.62 ;
        RECT  0.68 2.34 0.84 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.12 0.80 0.50 1.08 ;
        RECT  1.84 1.90 2.12 2.18 ;
        RECT  0.12 2.02 2.12 2.18 ;
        RECT  0.12 0.80 0.28 2.62 ;
        RECT  1.14 2.02 1.30 2.62 ;
        RECT  0.10 2.34 0.38 2.62 ;
        RECT  1.14 2.34 1.42 2.62 ;
        RECT  2.02 0.80 2.44 1.08 ;
        RECT  2.28 1.46 2.78 1.74 ;
        RECT  2.28 0.80 2.44 2.62 ;
        RECT  2.18 2.34 2.46 2.62 ;
        RECT  3.12 0.66 3.40 0.94 ;
        RECT  3.12 0.66 3.28 1.23 ;
        RECT  2.94 1.07 3.28 1.23 ;
        RECT  3.82 1.46 4.10 1.74 ;
        RECT  3.82 1.46 3.98 2.13 ;
        RECT  2.94 1.97 3.98 2.13 ;
        RECT  2.94 1.07 3.10 2.66 ;
        RECT  2.74 2.26 3.10 2.66 ;
    END
END AND3OR2SP2V1_0

MACRO AND3OR2SP1V1_0
    CLASS CORE ;
    FOREIGN AND3OR2SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.44 1.32 0.72 1.74 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.92 1.32 1.20 1.74 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.40 1.46 1.94 1.74 ;
        END
    END IN3
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 8.15  LAYER ME1  ;
        ANTENNADIFFAREA 3.47  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        ANTENNAMAXAREACAR 40.43  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.16 2.29 4.68 2.45 ;
        RECT  4.52 0.76 4.68 2.45 ;
        RECT  4.16 0.76 4.68 0.92 ;
        RECT  4.16 2.29 4.44 2.57 ;
        RECT  4.16 0.64 4.44 0.92 ;
        END
    END OUT
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.26 1.39 3.54 1.81 ;
        END
    END IN4
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.80 0.28 ;
        RECT  4.34 -0.28 4.62 0.32 ;
        RECT  3.64 0.64 3.92 0.92 ;
        RECT  3.70 -0.28 3.86 0.92 ;
        RECT  2.60 0.64 2.88 0.92 ;
        RECT  2.66 -0.28 2.82 0.92 ;
        RECT  1.50 0.80 1.78 1.08 ;
        RECT  1.54 -0.28 1.70 1.08 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.80 3.48 ;
        RECT  4.34 2.88 4.62 3.48 ;
        RECT  3.64 2.29 3.92 2.57 ;
        RECT  3.70 2.29 3.86 3.48 ;
        RECT  1.66 2.34 1.94 2.62 ;
        RECT  1.72 2.34 1.88 3.48 ;
        RECT  0.62 2.34 0.90 2.62 ;
        RECT  0.68 2.34 0.84 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.12 0.80 0.50 1.08 ;
        RECT  1.84 1.90 2.12 2.18 ;
        RECT  0.12 2.02 2.12 2.18 ;
        RECT  0.12 0.80 0.28 2.62 ;
        RECT  1.14 2.02 1.30 2.62 ;
        RECT  0.10 2.34 0.38 2.62 ;
        RECT  1.14 2.34 1.42 2.62 ;
        RECT  2.02 0.80 2.44 1.08 ;
        RECT  2.28 1.46 2.78 1.74 ;
        RECT  2.28 0.80 2.44 2.62 ;
        RECT  2.18 2.34 2.46 2.62 ;
        RECT  3.12 0.64 3.40 0.92 ;
        RECT  3.12 0.64 3.28 1.23 ;
        RECT  2.94 1.07 3.28 1.23 ;
        RECT  3.82 1.85 4.10 2.13 ;
        RECT  2.94 1.97 4.10 2.13 ;
        RECT  2.94 1.07 3.10 2.57 ;
        RECT  2.74 2.29 3.10 2.57 ;
    END
END AND3OR2SP1V1_0

MACRO AND3NOR2SP8V1_0
    CLASS CORE ;
    FOREIGN AND3NOR2SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 13.61  LAYER ME1  ;
        ANTENNADIFFAREA 7.87  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.64  LAYER ME1  ;
        ANTENNAMAXAREACAR 21.15  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.30 2.00 6.58 2.28 ;
        RECT  3.18 1.04 6.58 1.20 ;
        RECT  6.30 0.60 6.58 1.20 ;
        RECT  5.26 2.00 6.58 2.16 ;
        RECT  5.26 2.00 5.54 2.28 ;
        RECT  5.26 0.60 5.54 1.20 ;
        RECT  5.32 0.60 5.48 2.28 ;
        RECT  4.22 0.60 4.50 1.20 ;
        RECT  3.18 0.60 3.46 1.20 ;
        END
    END OUT
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.58  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.06 1.44 6.34 1.84 ;
        END
    END IN4
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.40 1.46 1.94 1.74 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.92 1.32 1.20 1.74 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.44 1.32 0.72 1.74 ;
        END
    END IN1
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 7.20 0.28 ;
        RECT  6.82 0.60 7.10 1.20 ;
        RECT  6.88 -0.28 7.04 1.20 ;
        RECT  6.74 -0.28 7.04 0.32 ;
        RECT  5.78 0.60 6.06 0.88 ;
        RECT  5.84 -0.28 6.00 0.88 ;
        RECT  4.74 0.60 5.02 0.88 ;
        RECT  4.80 -0.28 4.96 0.88 ;
        RECT  3.70 0.60 3.98 0.88 ;
        RECT  3.76 -0.28 3.92 0.88 ;
        RECT  2.66 0.60 2.94 1.20 ;
        RECT  2.72 -0.28 2.88 1.20 ;
        RECT  1.50 0.80 1.78 1.08 ;
        RECT  1.54 -0.28 1.70 1.08 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 7.20 3.48 ;
        RECT  6.74 2.88 7.02 3.48 ;
        RECT  4.22 2.32 4.50 2.60 ;
        RECT  4.28 2.32 4.44 3.48 ;
        RECT  3.18 2.32 3.46 2.60 ;
        RECT  3.24 2.32 3.40 3.48 ;
        RECT  1.66 2.34 1.94 2.62 ;
        RECT  1.72 2.34 1.88 3.48 ;
        RECT  0.62 2.34 0.90 2.62 ;
        RECT  0.68 2.34 0.84 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.12 0.80 0.50 1.08 ;
        RECT  1.80 1.90 2.08 2.18 ;
        RECT  0.12 2.02 2.08 2.18 ;
        RECT  0.12 0.80 0.28 2.62 ;
        RECT  1.14 2.02 1.30 2.62 ;
        RECT  0.10 2.34 0.38 2.62 ;
        RECT  1.14 2.34 1.42 2.62 ;
        RECT  2.02 0.80 2.40 1.08 ;
        RECT  2.24 1.52 3.10 1.68 ;
        RECT  2.82 1.46 3.10 1.74 ;
        RECT  2.24 0.80 2.40 2.62 ;
        RECT  2.18 2.34 2.46 2.62 ;
        RECT  2.66 2.00 5.02 2.16 ;
        RECT  4.74 2.00 5.02 2.60 ;
        RECT  5.78 2.32 6.06 2.60 ;
        RECT  2.66 2.00 2.94 2.60 ;
        RECT  3.70 2.00 3.98 2.60 ;
        RECT  6.82 2.00 7.10 2.60 ;
        RECT  4.74 2.44 7.10 2.60 ;
    END
END AND3NOR2SP8V1_0

MACRO AND3NOR2SP4V1_0
    CLASS CORE ;
    FOREIGN AND3NOR2SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.44 1.32 0.72 1.74 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.92 1.32 1.20 1.74 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.40 1.46 1.94 1.74 ;
        END
    END IN3
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.29  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.46 1.44 4.74 1.85 ;
        END
    END IN4
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 9.73  LAYER ME1  ;
        ANTENNADIFFAREA 5.07  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.36  LAYER ME1  ;
        ANTENNAMAXAREACAR 27.40  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.14 2.01 4.50 2.29 ;
        RECT  3.18 1.04 4.50 1.20 ;
        RECT  4.22 0.60 4.50 1.20 ;
        RECT  4.14 1.04 4.30 2.29 ;
        RECT  4.12 1.52 4.30 1.68 ;
        RECT  3.18 0.60 3.46 1.20 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 5.20 3.48 ;
        RECT  4.74 2.88 5.02 3.48 ;
        RECT  3.18 2.33 3.46 2.61 ;
        RECT  3.24 2.33 3.40 3.48 ;
        RECT  1.66 2.34 1.94 2.62 ;
        RECT  1.72 2.34 1.88 3.48 ;
        RECT  0.62 2.34 0.90 2.62 ;
        RECT  0.68 2.34 0.84 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 5.20 0.28 ;
        RECT  4.74 0.60 5.02 1.20 ;
        RECT  4.74 -0.28 5.02 0.32 ;
        RECT  4.80 -0.28 4.96 1.20 ;
        RECT  3.70 0.60 3.98 0.88 ;
        RECT  3.76 -0.28 3.92 0.88 ;
        RECT  2.66 0.60 2.94 1.20 ;
        RECT  2.72 -0.28 2.88 1.20 ;
        RECT  1.50 0.80 1.78 1.08 ;
        RECT  1.54 -0.28 1.70 1.08 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.12 0.80 0.50 1.08 ;
        RECT  1.80 1.90 2.08 2.18 ;
        RECT  0.12 2.02 2.08 2.18 ;
        RECT  0.12 0.80 0.28 2.62 ;
        RECT  1.14 2.02 1.30 2.62 ;
        RECT  0.10 2.34 0.38 2.62 ;
        RECT  1.14 2.34 1.42 2.62 ;
        RECT  2.02 0.80 2.40 1.08 ;
        RECT  2.24 1.52 3.10 1.68 ;
        RECT  2.82 1.46 3.10 1.74 ;
        RECT  2.24 0.80 2.40 2.62 ;
        RECT  2.18 2.34 2.46 2.62 ;
        RECT  2.66 2.01 3.98 2.17 ;
        RECT  3.70 2.01 3.98 2.61 ;
        RECT  2.66 2.01 2.94 2.61 ;
        RECT  4.74 2.01 5.02 2.61 ;
        RECT  3.70 2.45 5.02 2.61 ;
    END
END AND3NOR2SP4V1_0

MACRO AND3NOR2SP2V1_0
    CLASS CORE ;
    FOREIGN AND3NOR2SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 7.44  LAYER ME1  ;
        ANTENNADIFFAREA 3.71  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.21  LAYER ME1  ;
        ANTENNAMAXAREACAR 35.23  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.55 2.01 3.92 2.61 ;
        RECT  3.76 1.12 3.92 2.61 ;
        RECT  3.08 1.12 3.92 1.28 ;
        RECT  3.08 0.60 3.36 1.28 ;
        END
    END OUT
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.14  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.26 1.44 3.60 1.85 ;
        END
    END IN4
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.40 1.46 1.94 1.74 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.92 1.32 1.20 1.74 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.44 1.32 0.72 1.74 ;
        END
    END IN1
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.00 0.28 ;
        RECT  3.60 0.60 3.88 0.88 ;
        RECT  3.66 -0.28 3.82 0.88 ;
        RECT  3.54 -0.28 3.82 0.32 ;
        RECT  2.56 0.60 2.84 1.20 ;
        RECT  2.62 -0.28 2.78 1.20 ;
        RECT  1.50 0.80 1.78 1.08 ;
        RECT  1.54 -0.28 1.70 1.08 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.00 3.48 ;
        RECT  3.54 2.88 3.82 3.48 ;
        RECT  2.66 2.01 2.94 2.61 ;
        RECT  2.72 2.01 2.88 3.48 ;
        RECT  1.66 2.34 1.94 2.62 ;
        RECT  1.72 2.34 1.88 3.48 ;
        RECT  0.62 2.34 0.90 2.62 ;
        RECT  0.68 2.34 0.84 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.12 0.80 0.50 1.08 ;
        RECT  1.80 1.90 2.08 2.18 ;
        RECT  0.12 2.02 2.08 2.18 ;
        RECT  0.12 0.80 0.28 2.62 ;
        RECT  1.14 2.02 1.30 2.62 ;
        RECT  0.10 2.34 0.38 2.62 ;
        RECT  1.14 2.34 1.42 2.62 ;
        RECT  2.02 0.80 2.40 1.08 ;
        RECT  2.24 1.52 3.10 1.68 ;
        RECT  2.82 1.46 3.10 1.74 ;
        RECT  2.24 0.80 2.40 2.62 ;
        RECT  2.18 2.34 2.46 2.62 ;
    END
END AND3NOR2SP2V1_0

MACRO AND3NOR2SP1V1_0
    CLASS CORE ;
    FOREIGN AND3NOR2SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.44 1.32 0.72 1.74 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.92 1.32 1.20 1.74 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.40 1.46 1.94 1.74 ;
        END
    END IN3
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 6.70  LAYER ME1  ;
        ANTENNADIFFAREA 3.06  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        ANTENNAMAXAREACAR 49.86  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.55 2.02 3.92 2.30 ;
        RECT  3.76 1.12 3.92 2.30 ;
        RECT  3.21 1.12 3.92 1.28 ;
        RECT  3.21 0.63 3.37 1.28 ;
        RECT  3.09 0.63 3.37 0.91 ;
        END
    END OUT
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.26 1.44 3.60 1.86 ;
        END
    END IN4
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.00 0.28 ;
        RECT  3.61 0.63 3.89 0.91 ;
        RECT  3.67 -0.28 3.83 0.91 ;
        RECT  3.54 -0.28 3.83 0.32 ;
        RECT  2.57 0.63 2.85 0.91 ;
        RECT  2.63 -0.28 2.79 0.91 ;
        RECT  1.50 0.80 1.78 1.08 ;
        RECT  1.54 -0.28 1.70 1.08 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.00 3.48 ;
        RECT  3.54 2.88 3.82 3.48 ;
        RECT  2.66 2.02 2.94 2.30 ;
        RECT  2.72 2.02 2.88 3.48 ;
        RECT  1.66 2.34 1.94 2.62 ;
        RECT  1.72 2.34 1.88 3.48 ;
        RECT  0.62 2.34 0.90 2.62 ;
        RECT  0.68 2.34 0.84 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.12 0.80 0.50 1.08 ;
        RECT  1.80 1.90 2.08 2.18 ;
        RECT  0.12 2.02 2.08 2.18 ;
        RECT  0.12 0.80 0.28 2.62 ;
        RECT  1.14 2.02 1.30 2.62 ;
        RECT  0.10 2.34 0.38 2.62 ;
        RECT  1.14 2.34 1.42 2.62 ;
        RECT  2.02 0.80 2.40 1.08 ;
        RECT  2.24 1.52 3.10 1.68 ;
        RECT  2.82 1.46 3.10 1.74 ;
        RECT  2.24 0.80 2.40 2.62 ;
        RECT  2.18 2.34 2.46 2.62 ;
    END
END AND3NOR2SP1V1_0

MACRO AND3I2SP8V1_0
    CLASS CORE ;
    FOREIGN AND3I2SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 11.45  LAYER ME1  ;
        ANTENNADIFFAREA 6.40  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.92  LAYER ME1  ;
        ANTENNAMAXAREACAR 12.49  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.92 2.00 5.20 2.60 ;
        RECT  4.92 0.64 5.08 2.60 ;
        RECT  3.88 1.52 5.08 1.68 ;
        RECT  4.72 0.64 5.08 1.24 ;
        RECT  3.88 2.00 4.16 2.28 ;
        RECT  3.88 0.64 4.04 2.28 ;
        RECT  3.68 0.64 4.04 1.24 ;
        END
    END OUT
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.86 1.42 3.22 1.77 ;
        END
    END IN3
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.90 1.76 1.18 2.18 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.46 1.40 0.74 1.82 ;
        END
    END IN2
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 6.00 0.28 ;
        RECT  5.30 -0.28 5.82 0.32 ;
        RECT  5.24 0.64 5.52 1.24 ;
        RECT  5.30 -0.28 5.46 1.24 ;
        RECT  4.20 0.64 4.48 1.24 ;
        RECT  4.26 -0.28 4.42 1.24 ;
        RECT  3.16 0.64 3.44 1.24 ;
        RECT  3.22 -0.28 3.38 1.24 ;
        RECT  0.76 0.96 1.04 1.24 ;
        RECT  0.82 -0.28 0.98 1.24 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 6.00 3.48 ;
        RECT  5.50 2.88 5.82 3.48 ;
        RECT  5.44 2.00 5.72 2.60 ;
        RECT  5.50 2.00 5.66 3.48 ;
        RECT  4.40 2.00 4.68 2.60 ;
        RECT  4.46 2.00 4.62 3.48 ;
        RECT  3.32 2.48 3.60 2.76 ;
        RECT  3.38 2.48 3.54 3.48 ;
        RECT  2.28 2.48 2.56 2.76 ;
        RECT  2.34 2.48 2.50 3.48 ;
        RECT  0.76 2.34 1.04 2.62 ;
        RECT  0.82 2.34 0.98 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.44 0.38 0.72 ;
        RECT  0.14 0.96 0.52 1.24 ;
        RECT  0.14 0.44 0.30 2.62 ;
        RECT  0.14 2.34 0.52 2.62 ;
        RECT  1.28 0.96 1.56 1.24 ;
        RECT  1.34 1.46 2.10 1.62 ;
        RECT  1.82 1.42 2.10 1.70 ;
        RECT  1.34 0.96 1.50 2.62 ;
        RECT  1.28 2.34 1.56 2.62 ;
        RECT  1.88 0.68 2.42 1.24 ;
        RECT  3.42 1.44 3.70 1.72 ;
        RECT  2.26 0.68 2.42 2.16 ;
        RECT  3.42 1.44 3.58 2.16 ;
        RECT  1.78 2.00 3.58 2.16 ;
        RECT  1.78 2.00 1.94 2.60 ;
        RECT  2.80 2.00 2.96 2.60 ;
        RECT  1.76 2.32 2.04 2.60 ;
        RECT  2.80 2.32 3.08 2.60 ;
    END
END AND3I2SP8V1_0

MACRO AND3I2SP4V1_0
    CLASS CORE ;
    FOREIGN AND3I2SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.46 1.40 0.74 1.82 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.90 1.76 1.18 2.18 ;
        END
    END IN1
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.86 1.42 3.22 1.77 ;
        END
    END IN3
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 8.59  LAYER ME1  ;
        ANTENNADIFFAREA 4.82  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER ME1  ;
        ANTENNAMAXAREACAR 13.66  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.88 1.52 4.28 1.68 ;
        RECT  3.88 2.00 4.16 2.28 ;
        RECT  3.88 0.64 4.04 2.28 ;
        RECT  3.68 0.64 4.04 1.24 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.80 3.48 ;
        RECT  4.40 2.00 4.68 2.60 ;
        RECT  4.34 2.88 4.62 3.48 ;
        RECT  4.46 2.00 4.62 3.48 ;
        RECT  3.32 2.48 3.60 2.76 ;
        RECT  3.38 2.48 3.54 3.48 ;
        RECT  2.28 2.48 2.56 2.76 ;
        RECT  2.34 2.48 2.50 3.48 ;
        RECT  0.76 2.34 1.04 2.62 ;
        RECT  0.82 2.34 0.98 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.80 0.28 ;
        RECT  4.26 -0.28 4.62 0.32 ;
        RECT  4.20 0.64 4.48 1.24 ;
        RECT  4.26 -0.28 4.42 1.24 ;
        RECT  3.16 0.64 3.44 1.24 ;
        RECT  3.22 -0.28 3.38 1.24 ;
        RECT  0.76 0.96 1.04 1.24 ;
        RECT  0.82 -0.28 0.98 1.24 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.44 0.38 0.72 ;
        RECT  0.14 0.96 0.52 1.24 ;
        RECT  0.14 0.44 0.30 2.62 ;
        RECT  0.14 2.34 0.52 2.62 ;
        RECT  1.28 0.96 1.56 1.24 ;
        RECT  1.34 1.46 2.10 1.62 ;
        RECT  1.82 1.42 2.10 1.70 ;
        RECT  1.34 0.96 1.50 2.62 ;
        RECT  1.28 2.34 1.56 2.62 ;
        RECT  1.88 0.68 2.42 1.24 ;
        RECT  3.42 1.44 3.70 1.72 ;
        RECT  2.26 0.68 2.42 2.16 ;
        RECT  3.42 1.44 3.58 2.16 ;
        RECT  1.78 2.00 3.58 2.16 ;
        RECT  1.78 2.00 1.94 2.60 ;
        RECT  2.80 2.00 2.96 2.60 ;
        RECT  1.76 2.32 2.04 2.60 ;
        RECT  2.80 2.32 3.08 2.60 ;
    END
END AND3I2SP4V1_0

MACRO AND3I2SP2V1_0
    CLASS CORE ;
    FOREIGN AND3I2SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 8.24  LAYER ME1  ;
        ANTENNADIFFAREA 4.08  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.35  LAYER ME1  ;
        ANTENNAMAXAREACAR 23.84  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.88 2.06 4.28 2.34 ;
        RECT  4.12 0.64 4.28 2.34 ;
        RECT  3.68 0.64 4.28 1.24 ;
        END
    END OUT
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.10  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.86 1.40 3.22 1.75 ;
        END
    END IN3
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.90 1.76 1.18 2.18 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.46 1.40 0.74 1.82 ;
        END
    END IN2
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.40 0.28 ;
        RECT  3.94 -0.28 4.22 0.32 ;
        RECT  3.16 0.64 3.44 1.24 ;
        RECT  3.22 -0.28 3.38 1.24 ;
        RECT  0.76 0.96 1.04 1.24 ;
        RECT  0.82 -0.28 0.98 1.24 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.40 3.48 ;
        RECT  3.94 2.88 4.22 3.48 ;
        RECT  3.32 2.48 3.60 2.76 ;
        RECT  3.38 2.48 3.54 3.48 ;
        RECT  2.28 2.48 2.56 2.76 ;
        RECT  2.34 2.48 2.50 3.48 ;
        RECT  0.76 2.34 1.04 2.62 ;
        RECT  0.82 2.34 0.98 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.44 0.38 0.72 ;
        RECT  0.14 0.96 0.52 1.24 ;
        RECT  0.14 0.44 0.30 2.62 ;
        RECT  0.14 2.34 0.52 2.62 ;
        RECT  1.28 0.96 1.56 1.24 ;
        RECT  1.34 1.46 2.10 1.62 ;
        RECT  1.82 1.40 2.10 1.68 ;
        RECT  1.34 0.96 1.50 2.62 ;
        RECT  1.28 2.34 1.56 2.62 ;
        RECT  1.88 0.84 2.42 1.24 ;
        RECT  3.50 1.44 3.78 1.72 ;
        RECT  2.26 0.84 2.42 2.16 ;
        RECT  3.50 1.44 3.66 2.16 ;
        RECT  1.78 2.00 3.66 2.16 ;
        RECT  1.78 2.00 1.94 2.60 ;
        RECT  2.80 2.00 2.96 2.60 ;
        RECT  1.76 2.32 2.04 2.60 ;
        RECT  2.80 2.32 3.08 2.60 ;
    END
END AND3I2SP2V1_0

MACRO AND3I2SP1V1_0
    CLASS CORE ;
    FOREIGN AND3I2SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 8.01  LAYER ME1  ;
        ANTENNADIFFAREA 3.23  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        ANTENNAMAXAREACAR 39.71  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.84 2.32 4.28 2.60 ;
        RECT  4.12 0.78 4.28 2.60 ;
        RECT  3.68 0.78 4.28 1.06 ;
        END
    END OUT
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.86 1.40 3.22 1.75 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.46 1.40 0.74 1.82 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.90 1.76 1.18 2.18 ;
        END
    END IN1
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.40 3.48 ;
        RECT  3.94 2.88 4.22 3.48 ;
        RECT  3.32 2.32 3.60 2.60 ;
        RECT  3.38 2.32 3.54 3.48 ;
        RECT  2.28 2.32 2.56 2.60 ;
        RECT  2.34 2.32 2.50 3.48 ;
        RECT  0.76 2.34 1.04 2.62 ;
        RECT  0.82 2.34 0.98 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.40 0.28 ;
        RECT  3.94 -0.28 4.22 0.32 ;
        RECT  3.16 0.78 3.44 1.06 ;
        RECT  3.22 -0.28 3.38 1.06 ;
        RECT  0.76 0.96 1.04 1.24 ;
        RECT  0.82 -0.28 0.98 1.24 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.44 0.38 0.72 ;
        RECT  0.14 0.96 0.52 1.24 ;
        RECT  0.14 0.44 0.30 2.62 ;
        RECT  0.14 2.34 0.52 2.62 ;
        RECT  1.28 0.96 1.56 1.24 ;
        RECT  1.34 1.46 2.10 1.62 ;
        RECT  1.82 1.40 2.10 1.68 ;
        RECT  1.34 0.96 1.50 2.62 ;
        RECT  1.28 2.34 1.56 2.62 ;
        RECT  1.88 0.78 2.42 1.06 ;
        RECT  2.26 0.78 2.42 2.16 ;
        RECT  3.50 1.88 3.78 2.16 ;
        RECT  1.78 2.00 3.78 2.16 ;
        RECT  1.78 2.00 1.94 2.60 ;
        RECT  2.80 2.00 2.96 2.60 ;
        RECT  1.76 2.32 2.04 2.60 ;
        RECT  2.80 2.32 3.08 2.60 ;
    END
END AND3I2SP1V1_0

MACRO AND3I1SP8V1_0
    CLASS CORE ;
    FOREIGN AND3I1SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.17  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.46 1.28 0.74 1.70 ;
        END
    END IN1
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 9.86  LAYER ME1  ;
        ANTENNADIFFAREA 6.85  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.74  LAYER ME1  ;
        ANTENNAMAXAREACAR 13.25  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.26 2.00 4.54 2.60 ;
        RECT  4.26 0.58 4.42 2.60 ;
        RECT  3.32 1.52 4.42 1.68 ;
        RECT  4.14 0.58 4.42 1.18 ;
        RECT  3.22 2.00 3.50 2.28 ;
        RECT  3.32 1.03 3.48 2.28 ;
        RECT  3.10 0.90 3.38 1.19 ;
        END
    END OUT
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.17  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.40 1.39 2.68 1.81 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.17  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.70 1.49 2.16 1.78 ;
        END
    END IN2
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 5.20 0.28 ;
        RECT  4.72 -0.28 5.02 0.32 ;
        RECT  4.66 0.58 4.94 1.18 ;
        RECT  4.72 -0.28 4.88 1.18 ;
        RECT  3.62 0.58 3.90 0.86 ;
        RECT  3.68 -0.28 3.84 0.86 ;
        RECT  2.54 0.46 2.82 1.16 ;
        RECT  2.60 -0.28 2.76 1.16 ;
        RECT  0.62 0.44 0.90 1.12 ;
        RECT  0.68 -0.28 0.84 1.12 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 5.20 3.48 ;
        RECT  4.78 2.00 5.06 2.60 ;
        RECT  4.74 2.88 5.02 3.48 ;
        RECT  4.84 2.00 5.00 3.48 ;
        RECT  3.74 2.00 4.02 2.60 ;
        RECT  3.80 2.00 3.96 3.48 ;
        RECT  2.66 2.48 2.94 2.76 ;
        RECT  2.72 2.48 2.88 3.48 ;
        RECT  1.62 2.48 1.90 2.76 ;
        RECT  1.68 2.48 1.84 3.48 ;
        RECT  0.62 2.48 0.90 2.76 ;
        RECT  0.68 2.48 0.84 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.44 0.38 1.12 ;
        RECT  0.94 1.54 1.22 1.82 ;
        RECT  0.14 0.44 0.30 2.34 ;
        RECT  0.14 1.90 1.10 2.06 ;
        RECT  0.94 1.54 1.10 2.06 ;
        RECT  0.10 2.06 0.38 2.34 ;
        RECT  1.26 0.46 1.54 1.16 ;
        RECT  2.88 1.46 3.16 1.74 ;
        RECT  1.38 0.46 1.54 2.13 ;
        RECT  2.88 1.46 3.04 2.13 ;
        RECT  1.30 1.97 3.04 2.13 ;
        RECT  1.30 1.97 1.46 2.56 ;
        RECT  2.20 1.97 2.36 2.60 ;
        RECT  1.10 2.28 1.46 2.56 ;
        RECT  2.14 2.32 2.42 2.60 ;
    END
END AND3I1SP8V1_0

MACRO AND3I1SP4V1_0
    CLASS CORE ;
    FOREIGN AND3I1SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.14  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.70 1.49 2.16 1.78 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.14  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.40 1.39 2.68 1.81 ;
        END
    END IN3
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 7.74  LAYER ME1  ;
        ANTENNADIFFAREA 4.94  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.43  LAYER ME1  ;
        ANTENNAMAXAREACAR 18.11  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.22 2.00 3.50 2.28 ;
        RECT  3.32 1.03 3.48 2.28 ;
        RECT  3.10 0.90 3.38 1.19 ;
        END
    END OUT
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.14  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.46 1.28 0.74 1.70 ;
        END
    END IN1
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.40 0.28 ;
        RECT  3.68 -0.28 4.22 0.32 ;
        RECT  3.62 0.58 3.90 0.86 ;
        RECT  3.68 -0.28 3.84 0.86 ;
        RECT  2.58 0.58 2.86 1.18 ;
        RECT  2.64 -0.28 2.80 1.18 ;
        RECT  0.62 0.44 0.90 1.02 ;
        RECT  0.68 -0.28 0.84 1.02 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.40 3.48 ;
        RECT  3.80 2.88 4.22 3.48 ;
        RECT  3.74 2.00 4.02 2.60 ;
        RECT  3.80 2.00 3.96 3.48 ;
        RECT  2.66 2.48 2.94 2.76 ;
        RECT  2.72 2.48 2.88 3.48 ;
        RECT  1.62 2.48 1.90 2.76 ;
        RECT  1.68 2.48 1.84 3.48 ;
        RECT  0.62 2.18 0.90 2.76 ;
        RECT  0.68 2.18 0.84 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.44 0.38 1.02 ;
        RECT  0.94 1.58 1.22 1.86 ;
        RECT  0.14 1.86 1.10 2.02 ;
        RECT  0.14 0.44 0.30 2.76 ;
        RECT  0.10 2.18 0.38 2.76 ;
        RECT  1.26 0.58 1.54 1.16 ;
        RECT  2.88 1.46 3.16 1.74 ;
        RECT  1.38 0.58 1.54 2.13 ;
        RECT  2.88 1.46 3.04 2.13 ;
        RECT  1.30 1.97 3.04 2.13 ;
        RECT  1.30 1.97 1.46 2.56 ;
        RECT  2.20 1.97 2.36 2.60 ;
        RECT  1.10 2.28 1.46 2.56 ;
        RECT  2.14 2.32 2.42 2.60 ;
    END
END AND3I1SP4V1_0

MACRO AND3I1SP2V1_0
    CLASS CORE ;
    FOREIGN AND3I1SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 6.33  LAYER ME1  ;
        ANTENNADIFFAREA 3.53  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.24  LAYER ME1  ;
        ANTENNAMAXAREACAR 26.36  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.22 2.00 3.50 2.28 ;
        RECT  3.32 0.63 3.48 2.28 ;
        RECT  3.10 0.63 3.48 1.23 ;
        END
    END OUT
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.10  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.40 1.39 2.68 1.81 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.10  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.66 1.46 2.11 1.75 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.10  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.46 1.78 0.74 2.20 ;
        END
    END IN1
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 3.60 3.48 ;
        RECT  3.14 2.88 3.42 3.48 ;
        RECT  2.66 2.32 2.94 2.60 ;
        RECT  2.72 2.32 2.88 3.48 ;
        RECT  1.62 2.32 1.90 2.60 ;
        RECT  1.68 2.32 1.84 3.48 ;
        RECT  0.62 2.36 0.90 2.76 ;
        RECT  0.68 2.36 0.84 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 3.60 0.28 ;
        RECT  3.14 -0.28 3.42 0.32 ;
        RECT  2.58 0.63 2.86 1.23 ;
        RECT  2.64 -0.28 2.80 1.23 ;
        RECT  0.62 0.68 0.90 1.08 ;
        RECT  0.67 -0.28 0.83 1.08 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.68 0.38 1.08 ;
        RECT  0.14 1.46 1.18 1.62 ;
        RECT  0.90 1.41 1.18 1.69 ;
        RECT  0.14 0.68 0.30 2.76 ;
        RECT  0.10 2.36 0.38 2.76 ;
        RECT  1.26 0.68 1.54 1.08 ;
        RECT  2.88 1.46 3.16 1.74 ;
        RECT  1.34 0.68 1.50 2.13 ;
        RECT  2.88 1.46 3.04 2.13 ;
        RECT  1.22 1.97 3.04 2.13 ;
        RECT  1.22 1.97 1.38 2.56 ;
        RECT  2.20 1.97 2.36 2.60 ;
        RECT  1.10 2.28 1.38 2.56 ;
        RECT  2.14 2.32 2.42 2.60 ;
    END
END AND3I1SP2V1_0

MACRO AND3I1SP1V1_0
    CLASS CORE ;
    FOREIGN AND3I1SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.46 1.76 0.74 2.18 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.92 1.40 2.28 1.75 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.44 1.40 2.74 1.75 ;
        END
    END IN3
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 6.20  LAYER ME1  ;
        ANTENNADIFFAREA 2.75  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        ANTENNAMAXAREACAR 46.11  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.18 2.32 3.48 2.60 ;
        RECT  3.32 0.78 3.48 2.60 ;
        RECT  3.02 0.78 3.48 1.06 ;
        END
    END OUT
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 3.60 0.28 ;
        RECT  3.14 -0.28 3.42 0.32 ;
        RECT  2.50 0.78 2.78 1.06 ;
        RECT  2.56 -0.28 2.72 1.06 ;
        RECT  0.62 0.80 0.90 1.08 ;
        RECT  0.68 -0.28 0.84 1.08 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 3.60 3.48 ;
        RECT  3.14 2.88 3.42 3.48 ;
        RECT  2.66 2.32 2.94 2.60 ;
        RECT  2.72 2.32 2.88 3.48 ;
        RECT  1.62 2.32 1.90 2.60 ;
        RECT  1.68 2.32 1.84 3.48 ;
        RECT  0.62 2.34 0.90 2.62 ;
        RECT  0.68 2.34 0.84 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.80 0.38 1.08 ;
        RECT  0.14 1.44 1.44 1.60 ;
        RECT  1.16 1.38 1.44 1.66 ;
        RECT  0.14 0.80 0.30 2.62 ;
        RECT  0.10 2.34 0.38 2.62 ;
        RECT  1.22 0.78 1.76 1.06 ;
        RECT  1.60 0.78 1.76 2.16 ;
        RECT  2.84 1.88 3.12 2.16 ;
        RECT  1.12 2.00 3.12 2.16 ;
        RECT  1.12 2.00 1.28 2.60 ;
        RECT  2.14 2.00 2.30 2.60 ;
        RECT  1.10 2.32 1.38 2.60 ;
        RECT  2.14 2.32 2.42 2.60 ;
    END
END AND3I1SP1V1_0

MACRO AND2SP8V1_0
    CLASS CORE ;
    FOREIGN AND2SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 7.89  LAYER ME1  ;
        ANTENNADIFFAREA 5.28  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.58  LAYER ME1  ;
        ANTENNAMAXAREACAR 13.70  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.74 1.97 3.02 2.57 ;
        RECT  2.74 0.54 3.02 1.14 ;
        RECT  2.74 0.54 2.90 2.57 ;
        RECT  1.82 1.52 2.90 1.68 ;
        RECT  1.70 1.97 1.98 2.57 ;
        RECT  1.82 0.71 1.98 2.57 ;
        RECT  1.70 0.71 1.98 0.99 ;
        END
    END OUT
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.17  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.17  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.00 3.48 ;
        RECT  3.32 2.88 3.82 3.48 ;
        RECT  3.26 1.97 3.54 2.57 ;
        RECT  3.32 1.97 3.48 3.48 ;
        RECT  2.22 1.97 2.50 2.57 ;
        RECT  2.28 1.97 2.44 3.48 ;
        RECT  1.14 1.97 1.42 2.67 ;
        RECT  1.20 1.97 1.36 3.48 ;
        RECT  0.10 1.97 0.38 2.67 ;
        RECT  0.16 1.97 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.00 0.28 ;
        RECT  3.32 -0.28 3.82 0.32 ;
        RECT  3.26 0.54 3.54 1.14 ;
        RECT  3.32 -0.28 3.48 1.14 ;
        RECT  2.22 0.54 2.50 1.14 ;
        RECT  2.28 -0.28 2.44 1.14 ;
        RECT  1.14 0.44 1.42 0.72 ;
        RECT  1.20 -0.28 1.36 0.72 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.24 0.44 0.70 1.14 ;
        RECT  0.54 1.07 1.54 1.23 ;
        RECT  1.38 1.07 1.54 1.74 ;
        RECT  1.38 1.46 1.66 1.74 ;
        RECT  0.54 0.44 0.70 2.55 ;
        RECT  0.62 1.97 0.90 2.67 ;
    END
END AND2SP8V1_0

MACRO AND2SP4V1_0
    CLASS CORE ;
    FOREIGN AND2SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 2.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.14  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.14  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 5.01  LAYER ME1  ;
        ANTENNADIFFAREA 3.22  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.29  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.39  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.82 1.52 2.28 1.68 ;
        RECT  1.70 1.97 1.98 2.57 ;
        RECT  1.82 0.71 1.98 2.57 ;
        RECT  1.70 0.71 1.98 0.99 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 2.80 3.48 ;
        RECT  2.28 2.88 2.62 3.48 ;
        RECT  2.22 1.97 2.50 2.57 ;
        RECT  2.28 1.97 2.44 3.48 ;
        RECT  1.18 1.97 1.46 2.57 ;
        RECT  1.24 1.97 1.40 3.48 ;
        RECT  0.10 1.97 0.38 2.55 ;
        RECT  0.16 1.97 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 2.80 0.28 ;
        RECT  2.28 -0.28 2.62 0.32 ;
        RECT  2.22 0.54 2.50 1.14 ;
        RECT  2.28 -0.28 2.44 1.14 ;
        RECT  1.18 0.54 1.46 0.82 ;
        RECT  1.24 -0.28 1.40 0.82 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.24 0.56 0.70 1.14 ;
        RECT  0.54 1.07 1.54 1.23 ;
        RECT  1.38 1.07 1.54 1.74 ;
        RECT  1.38 1.46 1.66 1.74 ;
        RECT  0.54 0.56 0.70 2.55 ;
        RECT  0.54 1.97 0.90 2.55 ;
    END
END AND2SP4V1_0

MACRO AND2SP2V1_0
    CLASS CORE ;
    FOREIGN AND2SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 2.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 3.97  LAYER ME1  ;
        ANTENNADIFFAREA 2.33  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.14  LAYER ME1  ;
        ANTENNAMAXAREACAR 27.56  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.70 1.97 2.28 2.13 ;
        RECT  2.12 0.83 2.28 2.13 ;
        RECT  1.70 0.83 2.28 0.99 ;
        RECT  1.70 1.97 1.98 2.57 ;
        RECT  1.70 0.71 1.98 0.99 ;
        END
    END OUT
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.10  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.10  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 2.40 0.28 ;
        RECT  1.94 -0.28 2.22 0.32 ;
        RECT  1.18 0.54 1.46 0.82 ;
        RECT  1.24 -0.28 1.40 0.82 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 2.40 3.48 ;
        RECT  1.94 2.88 2.22 3.48 ;
        RECT  1.18 1.97 1.46 2.57 ;
        RECT  1.24 1.97 1.40 3.48 ;
        RECT  0.10 1.97 0.38 2.37 ;
        RECT  0.16 1.97 0.32 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.24 0.74 0.70 1.14 ;
        RECT  0.54 1.07 1.56 1.23 ;
        RECT  1.40 1.07 1.56 1.74 ;
        RECT  1.40 1.46 1.68 1.74 ;
        RECT  0.54 0.74 0.70 2.37 ;
        RECT  0.54 1.97 0.90 2.37 ;
    END
END AND2SP2V1_0

MACRO AND2SP1V1_0
    CLASS CORE ;
    FOREIGN AND2SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 2.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 3.81  LAYER ME1  ;
        ANTENNADIFFAREA 1.69  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        ANTENNAMAXAREACAR 56.63  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.66 1.97 2.28 2.13 ;
        RECT  2.12 0.75 2.28 2.13 ;
        RECT  1.66 0.75 2.28 0.91 ;
        RECT  1.66 1.97 1.94 2.25 ;
        RECT  1.66 0.63 1.94 0.91 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 2.40 3.48 ;
        RECT  1.94 2.88 2.22 3.48 ;
        RECT  1.14 1.97 1.42 2.25 ;
        RECT  1.20 1.97 1.36 3.48 ;
        RECT  0.10 1.97 0.38 2.25 ;
        RECT  0.16 1.97 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 2.40 0.28 ;
        RECT  1.94 -0.28 2.22 0.32 ;
        RECT  1.14 0.63 1.42 0.91 ;
        RECT  1.20 -0.28 1.36 0.91 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.24 0.63 0.70 0.91 ;
        RECT  0.54 1.07 1.68 1.23 ;
        RECT  1.40 1.07 1.68 1.35 ;
        RECT  0.54 0.63 0.70 2.25 ;
        RECT  0.54 1.97 0.90 2.25 ;
    END
END AND2SP1V1_0

MACRO AND2OR3SP8V1_0
    CLASS CORE ;
    FOREIGN AND2OR3SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 12.18  LAYER ME1  ;
        ANTENNADIFFAREA 6.93  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.81  LAYER ME1  ;
        ANTENNAMAXAREACAR 15.02  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.24 0.56 5.52 1.16 ;
        RECT  5.09 2.06 5.40 2.66 ;
        RECT  5.24 0.56 5.40 2.66 ;
        RECT  4.32 1.52 5.40 1.68 ;
        RECT  4.32 0.72 4.48 1.86 ;
        RECT  4.05 2.06 4.33 2.66 ;
        RECT  4.17 1.70 4.33 2.66 ;
        RECT  4.20 0.72 4.48 1.00 ;
        END
    END OUT
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.17  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.30 1.39 3.62 1.81 ;
        END
    END IN3
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.17  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.86 1.39 3.14 1.81 ;
        END
    END IN4
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 6.40 0.28 ;
        RECT  5.82 -0.28 6.22 0.32 ;
        RECT  5.76 0.56 6.04 1.16 ;
        RECT  5.82 -0.28 5.98 1.16 ;
        RECT  4.72 0.56 5.00 1.16 ;
        RECT  4.78 -0.28 4.94 1.16 ;
        RECT  3.64 0.44 3.92 0.72 ;
        RECT  3.70 -0.28 3.86 0.72 ;
        RECT  2.60 0.44 2.88 0.72 ;
        RECT  2.66 -0.28 2.82 0.72 ;
        RECT  1.04 0.63 1.32 0.91 ;
        RECT  1.10 -0.28 1.26 0.91 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 6.40 3.48 ;
        RECT  5.67 2.88 6.22 3.48 ;
        RECT  5.61 2.06 5.89 2.66 ;
        RECT  5.67 2.06 5.83 3.48 ;
        RECT  4.57 2.06 4.85 2.66 ;
        RECT  4.63 2.06 4.79 3.48 ;
        RECT  3.49 2.06 3.77 2.76 ;
        RECT  3.55 2.06 3.71 3.48 ;
        RECT  1.14 1.97 1.42 2.25 ;
        RECT  1.20 1.97 1.36 3.48 ;
        RECT  0.10 1.97 0.38 2.25 ;
        RECT  0.16 1.97 0.32 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.14 0.63 0.70 0.91 ;
        RECT  0.54 1.07 1.60 1.23 ;
        RECT  1.32 1.07 1.60 1.35 ;
        RECT  0.54 0.63 0.70 2.25 ;
        RECT  0.54 1.97 0.90 2.25 ;
        RECT  1.56 0.63 1.92 0.91 ;
        RECT  1.76 1.45 2.38 1.61 ;
        RECT  2.10 1.39 2.38 1.67 ;
        RECT  1.76 0.63 1.92 2.25 ;
        RECT  1.66 1.97 1.94 2.25 ;
        RECT  3.12 0.51 3.40 0.79 ;
        RECT  2.08 0.56 2.36 0.84 ;
        RECT  2.20 0.56 2.36 1.23 ;
        RECT  3.18 0.51 3.34 1.23 ;
        RECT  2.20 1.07 4.02 1.23 ;
        RECT  3.86 1.07 4.02 1.54 ;
        RECT  3.86 1.26 4.14 1.54 ;
        RECT  2.54 1.07 2.70 2.76 ;
        RECT  2.21 2.06 2.70 2.76 ;
    END
END AND2OR3SP8V1_0

MACRO AND2OR3SP4V1_0
    CLASS CORE ;
    FOREIGN AND2OR3SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.14  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.86 1.39 3.14 1.81 ;
        END
    END IN4
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.14  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.30 1.39 3.62 1.81 ;
        END
    END IN3
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 9.75  LAYER ME1  ;
        ANTENNADIFFAREA 5.27  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER ME1  ;
        ANTENNAMAXAREACAR 19.72  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.32 1.52 4.68 1.68 ;
        RECT  4.32 0.72 4.48 1.86 ;
        RECT  4.05 2.06 4.33 2.66 ;
        RECT  4.17 1.70 4.33 2.66 ;
        RECT  4.20 0.72 4.48 1.00 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 5.20 3.48 ;
        RECT  4.63 2.88 5.02 3.48 ;
        RECT  4.57 2.06 4.85 2.66 ;
        RECT  4.63 2.06 4.79 3.48 ;
        RECT  3.53 2.06 3.81 2.66 ;
        RECT  3.59 2.06 3.75 3.48 ;
        RECT  1.14 1.97 1.42 2.25 ;
        RECT  1.20 1.97 1.36 3.48 ;
        RECT  0.10 1.97 0.38 2.25 ;
        RECT  0.16 1.97 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 5.20 0.28 ;
        RECT  4.74 -0.28 5.02 0.32 ;
        RECT  4.72 0.56 5.00 1.16 ;
        RECT  4.78 -0.28 4.94 1.16 ;
        RECT  3.68 0.56 3.96 0.84 ;
        RECT  3.74 -0.28 3.90 0.84 ;
        RECT  2.60 0.56 2.88 0.84 ;
        RECT  2.66 -0.28 2.82 0.84 ;
        RECT  1.04 0.63 1.32 0.91 ;
        RECT  1.10 -0.28 1.26 0.91 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.14 0.63 0.70 0.91 ;
        RECT  0.54 1.07 1.60 1.23 ;
        RECT  1.32 1.07 1.60 1.35 ;
        RECT  0.54 0.63 0.70 2.25 ;
        RECT  0.54 1.97 0.90 2.25 ;
        RECT  1.56 0.63 1.92 0.91 ;
        RECT  1.76 1.45 2.38 1.61 ;
        RECT  2.10 1.39 2.38 1.67 ;
        RECT  1.76 0.63 1.92 2.25 ;
        RECT  1.66 1.97 1.94 2.25 ;
        RECT  3.12 0.63 3.40 0.91 ;
        RECT  2.08 0.68 2.36 0.96 ;
        RECT  2.20 0.68 2.36 1.23 ;
        RECT  3.18 0.63 3.34 1.23 ;
        RECT  2.20 1.07 4.02 1.23 ;
        RECT  3.86 1.07 4.02 1.54 ;
        RECT  3.86 1.26 4.14 1.54 ;
        RECT  2.54 1.07 2.70 2.65 ;
        RECT  2.21 2.07 2.70 2.65 ;
    END
END AND2OR3SP4V1_0

MACRO AND2OR3SP2V1_0
    CLASS CORE ;
    FOREIGN AND2OR3SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 9.01  LAYER ME1  ;
        ANTENNADIFFAREA 4.27  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.31  LAYER ME1  ;
        ANTENNAMAXAREACAR 29.32  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.05 2.06 4.68 2.66 ;
        RECT  4.52 0.70 4.68 2.66 ;
        RECT  4.20 0.70 4.68 0.98 ;
        END
    END OUT
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.10  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.30 1.39 3.62 1.81 ;
        END
    END IN3
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.10  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.86 1.39 3.14 1.81 ;
        END
    END IN4
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.80 3.48 ;
        RECT  4.34 2.88 4.62 3.48 ;
        RECT  3.53 2.06 3.81 2.66 ;
        RECT  3.59 2.06 3.75 3.48 ;
        RECT  1.14 1.97 1.42 2.25 ;
        RECT  1.20 1.97 1.36 3.48 ;
        RECT  0.10 1.97 0.38 2.25 ;
        RECT  0.16 1.97 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.80 0.28 ;
        RECT  4.38 -0.28 4.66 0.32 ;
        RECT  3.68 0.54 3.96 0.82 ;
        RECT  3.74 -0.28 3.90 0.82 ;
        RECT  2.60 0.54 2.88 0.82 ;
        RECT  2.66 -0.28 2.82 0.82 ;
        RECT  1.04 0.63 1.32 0.91 ;
        RECT  1.10 -0.28 1.26 0.91 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.14 0.63 0.70 0.91 ;
        RECT  0.54 1.07 1.60 1.23 ;
        RECT  1.32 1.07 1.60 1.35 ;
        RECT  0.54 0.63 0.70 2.25 ;
        RECT  0.54 1.97 0.90 2.25 ;
        RECT  1.56 0.63 1.92 0.91 ;
        RECT  1.76 1.45 2.38 1.61 ;
        RECT  2.10 1.39 2.38 1.67 ;
        RECT  1.76 0.63 1.92 2.25 ;
        RECT  1.66 1.97 1.94 2.25 ;
        RECT  3.12 0.63 3.40 0.91 ;
        RECT  2.08 0.66 2.36 0.94 ;
        RECT  2.20 0.66 2.36 1.23 ;
        RECT  3.18 0.63 3.34 1.23 ;
        RECT  2.20 1.07 4.02 1.23 ;
        RECT  3.86 1.07 4.02 1.54 ;
        RECT  3.86 1.26 4.14 1.54 ;
        RECT  2.54 1.07 2.70 2.47 ;
        RECT  2.21 2.07 2.70 2.47 ;
    END
END AND2OR3SP2V1_0

MACRO AND2OR3SP1V1_0
    CLASS CORE ;
    FOREIGN AND2OR3SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 8.76  LAYER ME1  ;
        ANTENNADIFFAREA 3.89  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.23  LAYER ME1  ;
        ANTENNAMAXAREACAR 38.03  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.05 2.07 4.68 2.35 ;
        RECT  4.52 0.66 4.68 2.35 ;
        RECT  4.20 0.66 4.68 0.94 ;
        END
    END OUT
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.10  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.30 1.39 3.62 1.81 ;
        END
    END IN3
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.10  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.86 1.39 3.14 1.81 ;
        END
    END IN4
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.80 0.28 ;
        RECT  4.38 -0.28 4.66 0.32 ;
        RECT  3.64 0.54 3.92 0.82 ;
        RECT  3.70 -0.28 3.86 0.82 ;
        RECT  2.60 0.54 2.88 0.82 ;
        RECT  2.66 -0.28 2.82 0.82 ;
        RECT  1.04 0.63 1.32 0.91 ;
        RECT  1.10 -0.28 1.26 0.91 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.80 3.48 ;
        RECT  4.34 2.88 4.62 3.48 ;
        RECT  3.49 2.07 3.77 2.47 ;
        RECT  3.55 2.07 3.71 3.48 ;
        RECT  1.14 1.97 1.42 2.25 ;
        RECT  1.20 1.97 1.36 3.48 ;
        RECT  0.10 1.97 0.38 2.25 ;
        RECT  0.16 1.97 0.32 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.14 0.63 0.70 0.91 ;
        RECT  0.54 1.07 1.60 1.23 ;
        RECT  1.32 1.07 1.60 1.35 ;
        RECT  0.54 0.63 0.70 2.25 ;
        RECT  0.54 1.97 0.90 2.25 ;
        RECT  1.56 0.63 1.92 0.91 ;
        RECT  1.76 1.45 2.38 1.61 ;
        RECT  2.10 1.39 2.38 1.67 ;
        RECT  1.76 0.63 1.92 2.25 ;
        RECT  1.66 1.97 1.94 2.25 ;
        RECT  3.12 0.63 3.40 0.91 ;
        RECT  2.08 0.66 2.36 0.94 ;
        RECT  2.20 0.66 2.36 1.23 ;
        RECT  3.18 0.63 3.34 1.23 ;
        RECT  2.20 1.07 4.02 1.23 ;
        RECT  3.86 1.09 4.14 1.37 ;
        RECT  2.54 1.07 2.70 2.47 ;
        RECT  2.21 2.07 2.70 2.47 ;
    END
END AND2OR3SP1V1_0

MACRO AND2OR2SP8V1_0
    CLASS CORE ;
    FOREIGN AND2OR2SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 11.76  LAYER ME1  ;
        ANTENNADIFFAREA 6.32  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.81  LAYER ME1  ;
        ANTENNAMAXAREACAR 14.49  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.78 0.54 5.06 1.14 ;
        RECT  4.66 2.06 4.94 2.66 ;
        RECT  4.78 0.54 4.94 2.66 ;
        RECT  3.82 1.52 4.94 1.68 ;
        RECT  3.74 0.86 4.02 1.14 ;
        RECT  3.62 2.06 3.98 2.66 ;
        RECT  3.82 0.86 3.98 2.66 ;
        END
    END OUT
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.17  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.90 1.42 3.18 1.84 ;
        END
    END IN3
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 6.00 0.28 ;
        RECT  5.36 -0.28 5.82 0.32 ;
        RECT  5.30 0.54 5.58 1.14 ;
        RECT  5.36 -0.28 5.52 1.14 ;
        RECT  4.26 0.54 4.54 1.14 ;
        RECT  4.32 -0.28 4.48 1.14 ;
        RECT  3.18 0.44 3.46 0.72 ;
        RECT  3.24 -0.28 3.40 0.72 ;
        RECT  2.14 0.44 2.42 1.14 ;
        RECT  2.20 -0.28 2.36 1.14 ;
        RECT  1.14 0.63 1.42 0.91 ;
        RECT  1.20 -0.28 1.36 0.91 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 6.00 3.48 ;
        RECT  5.24 2.88 5.82 3.48 ;
        RECT  5.18 2.06 5.46 2.66 ;
        RECT  5.24 2.06 5.40 3.48 ;
        RECT  4.14 2.06 4.42 2.66 ;
        RECT  4.20 2.06 4.36 3.48 ;
        RECT  3.06 2.06 3.34 2.76 ;
        RECT  3.12 2.06 3.28 3.48 ;
        RECT  1.14 1.97 1.42 2.25 ;
        RECT  1.20 1.97 1.36 3.48 ;
        RECT  0.10 1.97 0.38 2.25 ;
        RECT  0.16 1.97 0.32 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.24 0.63 0.70 0.91 ;
        RECT  0.54 1.07 1.60 1.23 ;
        RECT  1.32 1.07 1.60 1.35 ;
        RECT  0.54 0.63 0.70 2.25 ;
        RECT  0.54 1.97 0.90 2.25 ;
        RECT  1.66 0.63 1.94 0.91 ;
        RECT  1.76 1.40 2.42 1.56 ;
        RECT  2.14 1.34 2.42 1.62 ;
        RECT  1.76 0.63 1.92 2.25 ;
        RECT  1.66 1.97 1.94 2.25 ;
        RECT  2.58 0.44 2.94 1.26 ;
        RECT  2.58 1.10 3.54 1.26 ;
        RECT  3.38 1.10 3.54 1.81 ;
        RECT  3.38 1.53 3.66 1.81 ;
        RECT  2.58 0.44 2.74 2.76 ;
        RECT  2.16 2.06 2.74 2.76 ;
    END
END AND2OR2SP8V1_0

MACRO AND2OR2SP4V1_0
    CLASS CORE ;
    FOREIGN AND2OR2SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.14  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.90 1.42 3.18 1.84 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 9.30  LAYER ME1  ;
        ANTENNADIFFAREA 4.77  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER ME1  ;
        ANTENNAMAXAREACAR 18.81  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.82 1.52 4.28 1.68 ;
        RECT  3.74 0.86 4.02 1.14 ;
        RECT  3.62 2.00 3.98 2.60 ;
        RECT  3.82 0.86 3.98 2.60 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.80 3.48 ;
        RECT  4.20 2.88 4.62 3.48 ;
        RECT  4.14 2.00 4.42 2.60 ;
        RECT  4.20 2.00 4.36 3.48 ;
        RECT  3.10 2.00 3.38 2.60 ;
        RECT  3.16 2.00 3.32 3.48 ;
        RECT  1.14 1.97 1.42 2.25 ;
        RECT  1.20 1.97 1.36 3.48 ;
        RECT  0.10 1.97 0.38 2.25 ;
        RECT  0.16 1.97 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.80 0.28 ;
        RECT  4.32 -0.28 4.62 0.32 ;
        RECT  4.26 0.54 4.54 1.14 ;
        RECT  4.32 -0.28 4.48 1.14 ;
        RECT  3.18 0.44 3.46 0.72 ;
        RECT  3.24 -0.28 3.40 0.72 ;
        RECT  2.14 0.44 2.42 1.02 ;
        RECT  2.20 -0.28 2.36 1.02 ;
        RECT  1.14 0.63 1.42 0.91 ;
        RECT  1.20 -0.28 1.36 0.91 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.24 0.63 0.70 0.91 ;
        RECT  0.54 1.07 1.60 1.23 ;
        RECT  1.32 1.07 1.60 1.35 ;
        RECT  0.54 0.63 0.70 2.25 ;
        RECT  0.54 1.97 0.90 2.25 ;
        RECT  1.66 0.63 1.94 0.91 ;
        RECT  1.76 1.40 2.42 1.56 ;
        RECT  2.14 1.34 2.42 1.62 ;
        RECT  1.76 0.63 1.92 2.25 ;
        RECT  1.66 1.97 1.94 2.25 ;
        RECT  2.58 0.44 2.94 1.18 ;
        RECT  2.58 1.02 3.54 1.18 ;
        RECT  3.38 1.02 3.54 1.81 ;
        RECT  3.38 1.53 3.66 1.81 ;
        RECT  2.58 0.44 2.74 2.58 ;
        RECT  2.16 2.00 2.74 2.58 ;
    END
END AND2OR2SP4V1_0

MACRO AND2OR2SP2V1_0
    CLASS CORE ;
    FOREIGN AND2OR2SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 8.26  LAYER ME1  ;
        ANTENNADIFFAREA 3.86  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.31  LAYER ME1  ;
        ANTENNAMAXAREACAR 26.89  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.60 2.00 4.28 2.16 ;
        RECT  4.12 0.98 4.28 2.16 ;
        RECT  3.74 0.98 4.28 1.14 ;
        RECT  3.74 0.86 4.02 1.14 ;
        RECT  3.60 2.00 3.88 2.60 ;
        END
    END OUT
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.10  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.90 1.42 3.18 1.84 ;
        END
    END IN3
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.40 0.28 ;
        RECT  3.94 -0.28 4.22 0.32 ;
        RECT  3.22 0.54 3.50 0.82 ;
        RECT  3.28 -0.28 3.44 0.82 ;
        RECT  2.14 0.54 2.42 0.94 ;
        RECT  2.20 -0.28 2.36 0.94 ;
        RECT  1.14 0.63 1.42 0.91 ;
        RECT  1.20 -0.28 1.36 0.91 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.40 3.48 ;
        RECT  3.94 2.88 4.22 3.48 ;
        RECT  3.08 2.00 3.36 2.60 ;
        RECT  3.14 2.00 3.30 3.48 ;
        RECT  1.14 1.97 1.42 2.25 ;
        RECT  1.20 1.97 1.36 3.48 ;
        RECT  0.10 1.97 0.38 2.25 ;
        RECT  0.16 1.97 0.32 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.24 0.63 0.70 0.91 ;
        RECT  0.54 1.07 1.60 1.23 ;
        RECT  1.32 1.07 1.60 1.35 ;
        RECT  0.54 0.63 0.70 2.25 ;
        RECT  0.54 1.97 0.90 2.25 ;
        RECT  1.66 0.63 1.94 0.91 ;
        RECT  1.76 1.40 2.42 1.56 ;
        RECT  2.14 1.34 2.42 1.62 ;
        RECT  1.76 0.63 1.92 2.25 ;
        RECT  1.66 1.97 1.94 2.25 ;
        RECT  2.58 0.54 2.94 0.94 ;
        RECT  2.58 1.10 3.56 1.26 ;
        RECT  3.40 1.10 3.56 1.81 ;
        RECT  3.40 1.53 3.68 1.81 ;
        RECT  2.58 0.54 2.74 2.40 ;
        RECT  2.14 2.00 2.74 2.40 ;
    END
END AND2OR2SP2V1_0

MACRO AND2OR2SP1V1_0
    CLASS CORE ;
    FOREIGN AND2OR2SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 7.50  LAYER ME1  ;
        ANTENNADIFFAREA 3.22  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        ANTENNAMAXAREACAR 37.21  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.70 1.97 4.28 2.13 ;
        RECT  4.12 0.74 4.28 2.13 ;
        RECT  3.70 0.74 4.28 0.90 ;
        RECT  3.70 1.97 3.98 2.25 ;
        RECT  3.70 0.62 3.98 0.90 ;
        END
    END OUT
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.90 1.06 3.18 1.48 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.40 0.28 ;
        RECT  3.94 -0.28 4.22 0.32 ;
        RECT  3.18 0.62 3.46 0.90 ;
        RECT  3.24 -0.28 3.40 0.90 ;
        RECT  2.14 0.62 2.42 0.90 ;
        RECT  2.20 -0.28 2.36 0.90 ;
        RECT  1.14 0.63 1.42 0.91 ;
        RECT  1.20 -0.28 1.36 0.91 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.40 3.48 ;
        RECT  3.94 2.88 4.22 3.48 ;
        RECT  3.18 1.97 3.46 2.25 ;
        RECT  3.24 1.97 3.40 3.48 ;
        RECT  1.14 1.97 1.42 2.25 ;
        RECT  1.20 1.97 1.36 3.48 ;
        RECT  0.10 1.97 0.38 2.25 ;
        RECT  0.16 1.97 0.32 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.24 0.63 0.70 0.91 ;
        RECT  0.54 1.07 1.60 1.23 ;
        RECT  1.32 1.07 1.60 1.35 ;
        RECT  0.54 0.63 0.70 2.25 ;
        RECT  0.54 1.97 0.90 2.25 ;
        RECT  1.66 0.63 1.94 0.91 ;
        RECT  1.76 1.40 2.42 1.56 ;
        RECT  2.14 1.34 2.42 1.62 ;
        RECT  1.76 0.63 1.92 2.25 ;
        RECT  1.66 1.97 1.94 2.25 ;
        RECT  2.58 0.62 2.94 0.90 ;
        RECT  3.36 1.53 3.64 1.81 ;
        RECT  2.58 1.65 3.64 1.81 ;
        RECT  2.58 0.62 2.74 2.25 ;
        RECT  2.28 1.97 2.74 2.25 ;
    END
END AND2OR2SP1V1_0

MACRO AND2NOR3SP8V1_0
    CLASS CORE ;
    FOREIGN AND2NOR3SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.32 1.46 2.74 1.74 ;
        END
    END IN4
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.28 1.62 1.70 ;
        END
    END IN3
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.28 0.38 1.70 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.28 1.14 1.70 ;
        END
    END IN2
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 14.39  LAYER ME1  ;
        ANTENNADIFFAREA 7.22  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.78  LAYER ME1  ;
        ANTENNAMAXAREACAR 18.51  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.38 1.85 6.66 2.45 ;
        RECT  6.38 0.64 6.66 1.24 ;
        RECT  6.38 0.64 6.54 2.45 ;
        RECT  5.46 1.53 6.54 1.69 ;
        RECT  5.34 1.85 5.62 2.45 ;
        RECT  5.46 0.64 5.62 2.45 ;
        RECT  5.34 0.64 5.62 1.24 ;
        END
    END OUT
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 7.60 0.28 ;
        RECT  6.96 -0.28 7.42 0.32 ;
        RECT  6.90 0.64 7.18 1.24 ;
        RECT  6.96 -0.28 7.12 1.24 ;
        RECT  5.86 0.64 6.14 1.24 ;
        RECT  5.92 -0.28 6.08 1.24 ;
        RECT  4.82 0.64 5.10 1.24 ;
        RECT  4.88 -0.28 5.04 1.24 ;
        RECT  2.78 0.68 3.06 0.96 ;
        RECT  2.84 -0.28 3.00 0.96 ;
        RECT  1.04 0.62 1.32 0.90 ;
        RECT  1.10 -0.28 1.26 0.90 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 7.60 3.48 ;
        RECT  6.96 2.88 7.42 3.48 ;
        RECT  6.90 1.85 7.18 2.45 ;
        RECT  6.96 1.85 7.12 3.48 ;
        RECT  5.86 1.85 6.14 2.45 ;
        RECT  5.92 1.85 6.08 3.48 ;
        RECT  4.82 1.85 5.10 2.45 ;
        RECT  4.88 1.85 5.04 3.48 ;
        RECT  3.82 2.24 4.10 2.52 ;
        RECT  3.88 2.24 4.04 3.48 ;
        RECT  2.78 2.24 3.06 2.52 ;
        RECT  2.84 2.24 3.00 3.48 ;
        RECT  1.14 2.62 1.42 3.48 ;
        RECT  0.10 1.86 0.38 2.14 ;
        RECT  0.16 1.86 0.32 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.14 0.62 0.60 0.90 ;
        RECT  0.54 0.63 0.70 2.14 ;
        RECT  0.54 1.86 0.90 2.14 ;
        RECT  0.74 1.86 0.90 2.46 ;
        RECT  0.74 2.30 1.88 2.46 ;
        RECT  1.72 2.30 1.88 2.76 ;
        RECT  1.72 2.48 2.00 2.76 ;
        RECT  1.56 0.62 1.94 0.90 ;
        RECT  1.78 1.06 2.09 1.34 ;
        RECT  1.78 0.62 1.94 2.14 ;
        RECT  1.66 1.86 1.94 2.14 ;
        RECT  2.26 0.68 2.54 0.96 ;
        RECT  2.38 0.68 2.54 1.30 ;
        RECT  2.38 1.14 4.16 1.30 ;
        RECT  3.88 1.14 4.16 1.42 ;
        RECT  2.90 1.14 3.06 2.08 ;
        RECT  2.38 1.92 3.06 2.08 ;
        RECT  2.38 1.92 2.54 2.52 ;
        RECT  2.26 2.24 2.54 2.52 ;
        RECT  4.06 0.68 4.34 0.96 ;
        RECT  4.34 1.47 5.28 1.63 ;
        RECT  5.00 1.41 5.28 1.69 ;
        RECT  3.42 1.92 4.50 2.08 ;
        RECT  4.34 0.80 4.50 2.52 ;
        RECT  3.42 1.92 3.58 2.52 ;
        RECT  3.30 2.24 3.58 2.52 ;
        RECT  4.34 2.24 4.62 2.52 ;
    END
END AND2NOR3SP8V1_0

MACRO AND2NOR3SP4V1_0
    CLASS CORE ;
    FOREIGN AND2NOR3SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.29  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.06 1.39 4.34 1.81 ;
        END
    END IN3
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.29  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.66 1.39 5.94 1.81 ;
        END
    END IN4
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 11.86  LAYER ME1  ;
        ANTENNADIFFAREA 6.82  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.36  LAYER ME1  ;
        ANTENNAMAXAREACAR 33.38  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.14 2.00 5.50 2.28 ;
        RECT  5.14 1.52 5.30 2.28 ;
        RECT  2.66 1.04 5.20 1.20 ;
        RECT  4.92 0.60 5.20 1.20 ;
        RECT  4.92 1.52 5.30 1.68 ;
        RECT  4.92 0.60 5.08 1.68 ;
        RECT  3.70 0.60 3.98 1.20 ;
        RECT  2.66 0.60 2.94 1.20 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 6.40 3.48 ;
        RECT  5.94 2.88 6.22 3.48 ;
        RECT  2.66 2.32 2.94 2.60 ;
        RECT  2.72 2.32 2.88 3.48 ;
        RECT  1.14 1.97 1.42 2.25 ;
        RECT  1.20 1.97 1.36 3.48 ;
        RECT  0.10 1.97 0.38 2.25 ;
        RECT  0.16 1.97 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 6.40 0.28 ;
        RECT  5.94 -0.28 6.22 0.32 ;
        RECT  5.44 0.60 5.72 1.20 ;
        RECT  5.50 -0.28 5.66 1.20 ;
        RECT  4.31 0.60 4.59 0.88 ;
        RECT  4.37 -0.28 4.53 0.88 ;
        RECT  3.18 0.60 3.46 0.88 ;
        RECT  3.24 -0.28 3.40 0.88 ;
        RECT  2.14 0.60 2.42 1.20 ;
        RECT  2.20 -0.28 2.36 1.20 ;
        RECT  1.04 0.63 1.32 0.91 ;
        RECT  1.10 -0.28 1.26 0.91 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.14 0.63 0.70 0.91 ;
        RECT  0.54 1.07 1.58 1.23 ;
        RECT  1.30 1.07 1.58 1.35 ;
        RECT  0.54 0.63 0.70 2.25 ;
        RECT  0.54 1.97 0.90 2.25 ;
        RECT  1.56 0.63 1.90 0.91 ;
        RECT  1.74 1.46 2.50 1.62 ;
        RECT  2.22 1.46 2.50 1.74 ;
        RECT  1.74 0.63 1.90 2.25 ;
        RECT  1.66 1.97 1.94 2.25 ;
        RECT  2.14 2.00 4.50 2.16 ;
        RECT  4.22 2.00 4.50 2.28 ;
        RECT  2.14 2.00 2.42 2.60 ;
        RECT  3.18 2.00 3.46 2.60 ;
        RECT  3.70 2.32 3.98 2.60 ;
        RECT  4.70 2.32 4.98 2.60 ;
        RECT  5.74 2.00 6.02 2.60 ;
        RECT  3.70 2.44 6.02 2.60 ;
    END
END AND2NOR3SP4V1_0

MACRO AND2NOR3SP2V1_0
    CLASS CORE ;
    FOREIGN AND2NOR3SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 7.48  LAYER ME1  ;
        ANTENNADIFFAREA 3.91  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.21  LAYER ME1  ;
        ANTENNAMAXAREACAR 35.40  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.58 1.04 3.90 1.20 ;
        RECT  3.62 0.60 3.90 1.20 ;
        RECT  3.48 2.06 3.88 2.66 ;
        RECT  3.72 0.60 3.88 2.66 ;
        RECT  2.58 0.60 2.86 1.20 ;
        END
    END OUT
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.14  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.26 1.44 3.54 1.86 ;
        END
    END IN4
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.14  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.78 1.38 3.10 1.80 ;
        END
    END IN3
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.00 3.48 ;
        RECT  3.54 2.88 3.82 3.48 ;
        RECT  2.20 2.06 2.48 2.66 ;
        RECT  2.26 2.06 2.42 3.48 ;
        RECT  1.14 1.97 1.42 2.25 ;
        RECT  1.20 1.97 1.36 3.48 ;
        RECT  0.10 1.97 0.38 2.25 ;
        RECT  0.16 1.97 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.00 0.28 ;
        RECT  3.54 -0.28 3.82 0.32 ;
        RECT  3.10 0.60 3.38 0.88 ;
        RECT  3.16 -0.28 3.32 0.88 ;
        RECT  2.06 0.60 2.34 1.20 ;
        RECT  2.12 -0.28 2.28 1.20 ;
        RECT  1.04 0.63 1.32 0.91 ;
        RECT  1.10 -0.28 1.26 0.91 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.14 0.63 0.70 0.91 ;
        RECT  0.54 1.07 1.58 1.23 ;
        RECT  1.30 1.07 1.58 1.35 ;
        RECT  0.54 0.63 0.70 2.25 ;
        RECT  0.54 1.97 0.90 2.25 ;
        RECT  1.56 0.63 1.90 0.91 ;
        RECT  1.74 1.46 2.50 1.62 ;
        RECT  2.22 1.46 2.50 1.74 ;
        RECT  1.74 0.63 1.90 2.25 ;
        RECT  1.66 1.97 1.94 2.25 ;
    END
END AND2NOR3SP2V1_0

MACRO AND2NOR3SP1V1_0
    CLASS CORE ;
    FOREIGN AND2NOR3SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 7.42  LAYER ME1  ;
        ANTENNADIFFAREA 3.63  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.23  LAYER ME1  ;
        ANTENNAMAXAREACAR 32.91  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.62 0.68 3.90 0.96 ;
        RECT  3.48 2.16 3.88 2.56 ;
        RECT  3.72 1.12 3.88 2.56 ;
        RECT  3.62 0.68 3.78 1.28 ;
        RECT  2.70 1.12 3.88 1.28 ;
        RECT  2.70 0.68 2.86 1.28 ;
        RECT  2.58 0.68 2.86 0.96 ;
        END
    END OUT
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.08  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.26 1.44 3.54 1.86 ;
        END
    END IN4
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.08  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.68 1.44 3.00 1.86 ;
        END
    END IN3
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.00 0.28 ;
        RECT  3.54 -0.28 3.82 0.32 ;
        RECT  3.10 0.68 3.38 0.96 ;
        RECT  3.16 -0.28 3.32 0.96 ;
        RECT  2.06 0.68 2.34 0.96 ;
        RECT  2.12 -0.28 2.28 0.96 ;
        RECT  1.06 0.63 1.34 0.91 ;
        RECT  1.12 -0.28 1.28 0.91 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.00 3.48 ;
        RECT  3.54 2.88 3.82 3.48 ;
        RECT  2.20 2.16 2.48 2.56 ;
        RECT  2.26 2.16 2.42 3.48 ;
        RECT  1.18 1.97 1.46 2.57 ;
        RECT  1.24 1.97 1.40 3.48 ;
        RECT  0.10 1.97 0.38 2.25 ;
        RECT  0.16 1.97 0.32 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.12 0.63 0.70 0.91 ;
        RECT  0.54 1.07 1.46 1.23 ;
        RECT  1.30 1.07 1.46 1.75 ;
        RECT  1.30 1.47 1.62 1.75 ;
        RECT  0.54 0.63 0.70 2.25 ;
        RECT  0.54 1.97 0.90 2.25 ;
        RECT  1.58 0.68 1.86 0.96 ;
        RECT  1.70 0.68 1.86 1.33 ;
        RECT  1.78 1.46 2.50 1.62 ;
        RECT  2.22 1.46 2.50 1.74 ;
        RECT  1.78 1.17 1.94 2.57 ;
        RECT  1.70 1.97 1.98 2.57 ;
    END
END AND2NOR3SP1V1_0

MACRO AND2NOR2SP8V1_0
    CLASS CORE ;
    FOREIGN AND2NOR2SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 12.98  LAYER ME1  ;
        ANTENNADIFFAREA 7.37  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.64  LAYER ME1  ;
        ANTENNAMAXAREACAR 20.19  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.78 2.00 6.06 2.28 ;
        RECT  2.66 1.07 6.06 1.23 ;
        RECT  5.78 0.63 6.06 1.23 ;
        RECT  4.74 2.00 6.06 2.16 ;
        RECT  5.32 1.07 5.48 2.16 ;
        RECT  4.74 2.00 5.02 2.28 ;
        RECT  4.74 0.63 5.02 1.23 ;
        RECT  3.70 0.63 3.98 1.23 ;
        RECT  2.66 0.63 2.94 1.23 ;
        END
    END OUT
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.58  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.06 1.40 6.34 1.80 ;
        END
    END IN3
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 6.80 0.28 ;
        RECT  6.34 -0.28 6.62 0.32 ;
        RECT  6.30 0.63 6.58 1.23 ;
        RECT  6.36 -0.28 6.52 1.23 ;
        RECT  5.26 0.63 5.54 0.91 ;
        RECT  5.32 -0.28 5.48 0.91 ;
        RECT  4.22 0.63 4.50 0.91 ;
        RECT  4.28 -0.28 4.44 0.91 ;
        RECT  3.18 0.63 3.46 0.91 ;
        RECT  3.22 -0.28 3.38 0.91 ;
        RECT  2.14 0.63 2.42 1.23 ;
        RECT  2.20 -0.28 2.36 1.23 ;
        RECT  1.14 0.63 1.42 0.91 ;
        RECT  1.20 -0.28 1.36 0.91 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 6.80 3.48 ;
        RECT  6.34 2.88 6.62 3.48 ;
        RECT  3.70 2.32 3.98 2.60 ;
        RECT  3.76 2.32 3.92 3.48 ;
        RECT  2.66 2.32 2.94 2.60 ;
        RECT  2.72 2.32 2.88 3.48 ;
        RECT  1.14 1.97 1.42 2.25 ;
        RECT  1.20 1.97 1.36 3.48 ;
        RECT  0.10 1.97 0.38 2.25 ;
        RECT  0.16 1.97 0.32 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.24 0.63 0.70 0.91 ;
        RECT  0.54 1.07 1.60 1.23 ;
        RECT  1.32 1.07 1.60 1.35 ;
        RECT  0.54 0.63 0.70 2.25 ;
        RECT  0.54 1.97 0.90 2.25 ;
        RECT  1.66 0.63 1.94 0.91 ;
        RECT  1.76 1.52 2.70 1.68 ;
        RECT  2.42 1.46 2.70 1.74 ;
        RECT  1.76 0.63 1.92 2.25 ;
        RECT  1.66 1.97 1.94 2.25 ;
        RECT  2.14 2.00 4.50 2.16 ;
        RECT  4.22 2.00 4.50 2.60 ;
        RECT  5.26 2.32 5.54 2.60 ;
        RECT  2.14 2.00 2.42 2.60 ;
        RECT  3.18 2.00 3.46 2.60 ;
        RECT  6.30 2.00 6.58 2.60 ;
        RECT  4.22 2.44 6.58 2.60 ;
    END
END AND2NOR2SP8V1_0

MACRO AND2NOR2SP4V1_0
    CLASS CORE ;
    FOREIGN AND2NOR2SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.29  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.06 1.40 4.34 1.80 ;
        END
    END IN3
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 9.08  LAYER ME1  ;
        ANTENNADIFFAREA 4.81  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.36  LAYER ME1  ;
        ANTENNAMAXAREACAR 25.56  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.70 2.00 3.98 2.28 ;
        RECT  2.66 1.07 3.98 1.23 ;
        RECT  3.70 0.63 3.98 1.23 ;
        RECT  3.72 0.63 3.88 2.28 ;
        RECT  2.66 0.63 2.94 1.23 ;
        END
    END OUT
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.80 0.28 ;
        RECT  4.28 -0.28 4.62 0.32 ;
        RECT  4.22 0.63 4.50 1.23 ;
        RECT  4.28 -0.28 4.44 1.23 ;
        RECT  3.18 0.63 3.46 0.91 ;
        RECT  3.22 -0.28 3.38 0.91 ;
        RECT  2.14 0.63 2.42 1.23 ;
        RECT  2.20 -0.28 2.36 1.23 ;
        RECT  1.14 0.63 1.42 0.91 ;
        RECT  1.20 -0.28 1.36 0.91 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.80 3.48 ;
        RECT  4.34 2.88 4.62 3.48 ;
        RECT  2.66 2.32 2.94 2.60 ;
        RECT  2.72 2.32 2.88 3.48 ;
        RECT  1.14 1.97 1.42 2.25 ;
        RECT  1.20 1.97 1.36 3.48 ;
        RECT  0.10 1.97 0.38 2.25 ;
        RECT  0.16 1.97 0.32 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.24 0.63 0.70 0.91 ;
        RECT  0.54 1.07 1.60 1.23 ;
        RECT  1.32 1.07 1.60 1.35 ;
        RECT  0.54 0.63 0.70 2.25 ;
        RECT  0.54 1.97 0.90 2.25 ;
        RECT  1.66 0.63 1.94 0.91 ;
        RECT  1.76 1.52 2.70 1.68 ;
        RECT  2.42 1.46 2.70 1.74 ;
        RECT  1.76 0.63 1.92 2.25 ;
        RECT  1.66 1.97 1.94 2.25 ;
        RECT  2.14 2.00 3.46 2.16 ;
        RECT  3.18 2.00 3.46 2.60 ;
        RECT  2.14 2.00 2.42 2.60 ;
        RECT  4.22 2.00 4.50 2.60 ;
        RECT  3.18 2.44 4.50 2.60 ;
    END
END AND2NOR2SP4V1_0

MACRO AND2NOR2SP2V1_0
    CLASS CORE ;
    FOREIGN AND2NOR2SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 6.77  LAYER ME1  ;
        ANTENNADIFFAREA 3.40  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.21  LAYER ME1  ;
        ANTENNAMAXAREACAR 32.05  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.36 1.12 3.52 2.18 ;
        RECT  3.13 2.02 3.41 2.62 ;
        RECT  2.66 1.12 3.52 1.28 ;
        RECT  2.66 0.63 2.94 1.28 ;
        END
    END OUT
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.14  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.90 1.44 3.18 1.86 ;
        END
    END IN3
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 3.60 3.48 ;
        RECT  3.14 2.88 3.42 3.48 ;
        RECT  2.23 2.02 2.51 2.62 ;
        RECT  2.29 2.02 2.45 3.48 ;
        RECT  1.14 1.97 1.42 2.25 ;
        RECT  1.20 1.97 1.36 3.48 ;
        RECT  0.10 1.97 0.38 2.25 ;
        RECT  0.16 1.97 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 3.60 0.28 ;
        RECT  3.18 0.63 3.46 0.91 ;
        RECT  3.14 -0.28 3.42 0.32 ;
        RECT  3.22 -0.28 3.38 0.91 ;
        RECT  2.14 0.63 2.42 1.23 ;
        RECT  2.20 -0.28 2.36 1.23 ;
        RECT  1.14 0.63 1.42 0.91 ;
        RECT  1.20 -0.28 1.36 0.91 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.24 0.63 0.70 0.91 ;
        RECT  0.54 1.07 1.60 1.23 ;
        RECT  1.32 1.07 1.60 1.35 ;
        RECT  0.54 0.63 0.70 2.25 ;
        RECT  0.54 1.97 0.90 2.25 ;
        RECT  1.66 0.63 1.94 0.91 ;
        RECT  1.76 1.52 2.70 1.68 ;
        RECT  2.42 1.46 2.70 1.74 ;
        RECT  1.76 0.63 1.92 2.25 ;
        RECT  1.66 1.97 1.94 2.25 ;
    END
END AND2NOR2SP2V1_0

MACRO AND2NOR2SP1V1_0
    CLASS CORE ;
    FOREIGN AND2NOR2SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.90 1.44 3.18 1.86 ;
        END
    END IN3
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 6.06  LAYER ME1  ;
        ANTENNADIFFAREA 2.75  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        ANTENNAMAXAREACAR 45.10  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.13 2.02 3.52 2.30 ;
        RECT  3.36 1.12 3.52 2.30 ;
        RECT  2.78 1.12 3.52 1.28 ;
        RECT  2.78 0.63 2.94 1.28 ;
        RECT  2.66 0.63 2.94 0.91 ;
        END
    END OUT
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.39 1.14 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 3.60 0.28 ;
        RECT  3.18 0.63 3.46 0.91 ;
        RECT  3.14 -0.28 3.42 0.32 ;
        RECT  3.22 -0.28 3.38 0.91 ;
        RECT  2.14 0.63 2.42 0.91 ;
        RECT  2.20 -0.28 2.36 0.91 ;
        RECT  1.14 0.63 1.42 0.91 ;
        RECT  1.20 -0.28 1.36 0.91 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 3.60 3.48 ;
        RECT  3.14 2.88 3.42 3.48 ;
        RECT  2.23 2.02 2.51 2.30 ;
        RECT  2.29 2.02 2.45 3.48 ;
        RECT  1.14 1.97 1.42 2.25 ;
        RECT  1.20 1.97 1.36 3.48 ;
        RECT  0.10 1.97 0.38 2.25 ;
        RECT  0.16 1.97 0.32 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.24 0.63 0.70 0.91 ;
        RECT  0.54 1.07 1.60 1.23 ;
        RECT  1.32 1.07 1.60 1.35 ;
        RECT  0.54 0.63 0.70 2.25 ;
        RECT  0.54 1.97 0.90 2.25 ;
        RECT  1.66 0.63 1.94 0.91 ;
        RECT  1.76 1.52 2.70 1.68 ;
        RECT  2.42 1.46 2.70 1.74 ;
        RECT  1.76 0.63 1.92 2.25 ;
        RECT  1.66 1.97 1.94 2.25 ;
    END
END AND2NOR2SP1V1_0

MACRO AND2I1SP8V1_0
    CLASS CORE ;
    FOREIGN AND2I1SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 9.91  LAYER ME1  ;
        ANTENNADIFFAREA 6.48  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.74  LAYER ME1  ;
        ANTENNAMAXAREACAR 13.32  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.74 1.97 4.02 2.57 ;
        RECT  3.74 0.60 4.02 1.20 ;
        RECT  3.74 0.60 3.90 2.57 ;
        RECT  2.90 1.52 3.90 1.68 ;
        RECT  2.70 1.97 3.06 2.57 ;
        RECT  2.90 0.73 3.06 2.57 ;
        RECT  2.70 0.73 3.06 1.01 ;
        END
    END OUT
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.17  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.95 1.46 2.28 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.17  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.80 0.28 ;
        RECT  4.32 -0.28 4.62 0.32 ;
        RECT  4.26 0.60 4.54 1.20 ;
        RECT  4.32 -0.28 4.48 1.20 ;
        RECT  3.22 0.60 3.50 1.20 ;
        RECT  3.28 -0.28 3.44 1.20 ;
        RECT  2.14 0.50 2.42 0.78 ;
        RECT  2.20 -0.28 2.36 0.78 ;
        RECT  0.10 0.53 0.38 1.23 ;
        RECT  0.16 -0.28 0.32 1.23 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.80 3.48 ;
        RECT  4.32 2.88 4.62 3.48 ;
        RECT  4.26 1.97 4.54 2.57 ;
        RECT  4.32 1.97 4.48 3.48 ;
        RECT  3.22 1.97 3.50 2.57 ;
        RECT  3.28 1.97 3.44 3.48 ;
        RECT  2.14 1.97 2.42 2.67 ;
        RECT  2.20 1.97 2.36 3.48 ;
        RECT  1.10 1.97 1.38 2.67 ;
        RECT  1.16 1.97 1.32 3.48 ;
        RECT  0.10 1.97 0.38 2.67 ;
        RECT  0.16 1.97 0.32 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.53 0.90 1.23 ;
        RECT  0.74 1.52 1.38 1.68 ;
        RECT  1.10 1.46 1.38 1.74 ;
        RECT  0.74 0.53 0.90 2.67 ;
        RECT  0.62 1.97 0.90 2.67 ;
        RECT  1.24 0.50 1.52 1.20 ;
        RECT  1.24 0.62 1.72 1.20 ;
        RECT  1.56 1.14 2.60 1.30 ;
        RECT  2.44 1.14 2.60 1.75 ;
        RECT  2.44 1.47 2.72 1.75 ;
        RECT  1.56 0.62 1.72 2.67 ;
        RECT  1.56 1.97 1.90 2.67 ;
    END
END AND2I1SP8V1_0

MACRO AND2I1SP4V1_0
    CLASS CORE ;
    FOREIGN AND2I1SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.14  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.14  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.95 1.46 2.28 1.81 ;
        END
    END IN2
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 6.90  LAYER ME1  ;
        ANTENNADIFFAREA 4.26  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.43  LAYER ME1  ;
        ANTENNAMAXAREACAR 16.16  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.90 1.52 3.08 1.68 ;
        RECT  2.70 1.97 3.06 2.57 ;
        RECT  2.90 0.73 3.06 2.57 ;
        RECT  2.70 0.73 3.06 1.01 ;
        END
    END OUT
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 3.60 0.28 ;
        RECT  3.22 0.60 3.50 1.20 ;
        RECT  3.28 -0.28 3.44 1.20 ;
        RECT  3.14 -0.28 3.44 0.32 ;
        RECT  2.18 0.60 2.46 0.88 ;
        RECT  2.24 -0.28 2.40 0.88 ;
        RECT  0.10 0.65 0.38 1.23 ;
        RECT  0.16 -0.28 0.32 1.23 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 3.60 3.48 ;
        RECT  3.22 1.97 3.50 2.57 ;
        RECT  3.14 2.88 3.44 3.48 ;
        RECT  3.28 1.97 3.44 3.48 ;
        RECT  2.18 1.97 2.46 2.57 ;
        RECT  2.24 1.97 2.40 3.48 ;
        RECT  1.10 1.97 1.38 2.55 ;
        RECT  1.16 1.97 1.32 3.48 ;
        RECT  0.10 1.97 0.38 2.55 ;
        RECT  0.16 1.97 0.32 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.65 0.90 1.23 ;
        RECT  0.74 1.52 1.38 1.68 ;
        RECT  1.10 1.46 1.38 1.74 ;
        RECT  0.74 0.65 0.90 2.55 ;
        RECT  0.62 1.97 0.90 2.55 ;
        RECT  1.24 0.62 1.72 1.20 ;
        RECT  1.56 1.14 2.60 1.30 ;
        RECT  2.44 1.14 2.60 1.75 ;
        RECT  2.44 1.47 2.72 1.75 ;
        RECT  1.56 0.62 1.72 2.55 ;
        RECT  1.56 1.97 1.90 2.55 ;
    END
END AND2I1SP4V1_0

MACRO AND2I1SP2V1_0
    CLASS CORE ;
    FOREIGN AND2I1SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 5.71  LAYER ME1  ;
        ANTENNADIFFAREA 3.13  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.24  LAYER ME1  ;
        ANTENNAMAXAREACAR 23.79  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.70 1.97 3.08 2.57 ;
        RECT  2.92 0.73 3.08 2.57 ;
        RECT  2.70 0.73 3.08 1.01 ;
        END
    END OUT
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.10  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.95 1.46 2.28 1.81 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.10  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 3.20 3.48 ;
        RECT  2.74 2.88 3.02 3.48 ;
        RECT  2.18 1.97 2.46 2.57 ;
        RECT  2.24 1.97 2.40 3.48 ;
        RECT  1.10 1.97 1.38 2.37 ;
        RECT  1.16 1.97 1.32 3.48 ;
        RECT  0.10 1.97 0.38 2.37 ;
        RECT  0.16 1.97 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 3.20 0.28 ;
        RECT  2.74 -0.28 3.02 0.32 ;
        RECT  2.18 0.54 2.46 0.82 ;
        RECT  2.24 -0.28 2.40 0.82 ;
        RECT  0.10 0.51 0.38 0.91 ;
        RECT  0.16 -0.28 0.32 0.91 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.51 0.90 0.91 ;
        RECT  0.74 1.52 1.38 1.68 ;
        RECT  1.10 1.46 1.38 1.74 ;
        RECT  0.74 0.51 0.90 2.37 ;
        RECT  0.62 1.97 0.90 2.37 ;
        RECT  1.24 0.74 1.72 1.14 ;
        RECT  1.56 1.14 2.60 1.30 ;
        RECT  2.44 1.14 2.60 1.75 ;
        RECT  2.44 1.47 2.72 1.75 ;
        RECT  1.56 0.74 1.72 2.37 ;
        RECT  1.56 1.97 1.90 2.37 ;
    END
END AND2I1SP2V1_0

MACRO AND2I1SP1V1_0
    CLASS CORE ;
    FOREIGN AND2I1SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 5.46  LAYER ME1  ;
        ANTENNADIFFAREA 2.33  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        ANTENNAMAXAREACAR 40.66  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.92 0.75 3.08 2.13 ;
        RECT  2.66 1.97 2.94 2.25 ;
        RECT  2.66 0.63 2.94 0.91 ;
        END
    END OUT
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.95 1.46 2.34 1.74 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.39 0.38 1.81 ;
        END
    END IN1
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 3.20 0.28 ;
        RECT  2.74 -0.28 3.02 0.32 ;
        RECT  2.14 0.63 2.42 0.91 ;
        RECT  2.20 -0.28 2.36 0.91 ;
        RECT  0.10 0.63 0.38 0.91 ;
        RECT  0.16 -0.28 0.32 0.91 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 3.20 3.48 ;
        RECT  2.74 2.88 3.02 3.48 ;
        RECT  2.14 1.97 2.42 2.25 ;
        RECT  2.20 1.97 2.36 3.48 ;
        RECT  1.10 1.97 1.38 2.25 ;
        RECT  1.16 1.97 1.32 3.48 ;
        RECT  0.10 1.97 0.38 2.25 ;
        RECT  0.16 1.97 0.32 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.62 0.63 0.90 0.91 ;
        RECT  0.74 1.52 1.38 1.68 ;
        RECT  1.10 1.46 1.38 1.74 ;
        RECT  0.74 0.63 0.90 2.25 ;
        RECT  0.62 1.97 0.90 2.25 ;
        RECT  1.24 0.63 1.72 0.91 ;
        RECT  1.56 1.07 2.74 1.23 ;
        RECT  2.46 1.07 2.74 1.35 ;
        RECT  1.56 0.63 1.72 2.25 ;
        RECT  1.56 1.97 1.90 2.25 ;
    END
END AND2I1SP1V1_0

MACRO AND23OR3SP8V1_0
    CLASS CORE ;
    FOREIGN AND23OR3SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 13.78  LAYER ME1  ;
        ANTENNADIFFAREA 7.59  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.76  LAYER ME1  ;
        ANTENNAMAXAREACAR 18.05  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.06 1.52 7.48 1.68 ;
        RECT  6.92 1.96 7.22 2.46 ;
        RECT  7.06 0.74 7.22 2.46 ;
        RECT  6.92 0.74 7.22 1.24 ;
        END
    END OUT
    PIN IN6
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.61 1.52 3.93 1.82 ;
        RECT  3.61 1.46 3.89 1.82 ;
        END
    END IN6
    PIN IN5
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.85 1.40 3.13 1.82 ;
        END
    END IN5
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.10 1.40 2.38 1.82 ;
        END
    END IN4
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.40 1.62 1.82 ;
        END
    END IN3
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.40 0.38 1.82 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.40 1.14 1.82 ;
        END
    END IN2
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 8.00 0.28 ;
        RECT  7.50 -0.28 7.82 0.32 ;
        RECT  7.44 0.74 7.72 1.24 ;
        RECT  7.50 -0.28 7.66 1.24 ;
        RECT  6.40 0.74 6.68 1.24 ;
        RECT  6.46 -0.28 6.62 1.24 ;
        RECT  3.85 0.68 4.13 0.96 ;
        RECT  3.91 -0.28 4.07 0.96 ;
        RECT  1.14 0.84 1.42 1.12 ;
        RECT  1.20 -0.28 1.36 1.12 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 8.00 3.48 ;
        RECT  7.50 2.88 7.82 3.48 ;
        RECT  7.44 1.96 7.72 2.46 ;
        RECT  7.50 1.96 7.66 3.48 ;
        RECT  6.40 1.96 6.68 2.46 ;
        RECT  6.46 1.96 6.62 3.48 ;
        RECT  4.88 2.24 5.16 2.52 ;
        RECT  4.95 2.24 5.11 3.48 ;
        RECT  3.84 2.24 4.12 2.52 ;
        RECT  3.90 2.24 4.06 3.48 ;
        RECT  2.76 1.98 3.04 2.26 ;
        RECT  2.82 1.98 2.98 3.48 ;
        RECT  1.14 1.98 1.42 2.26 ;
        RECT  1.20 1.98 1.36 3.48 ;
        RECT  0.10 1.98 0.38 2.26 ;
        RECT  0.16 1.98 0.32 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.44 0.38 0.72 ;
        RECT  0.22 0.44 0.38 1.12 ;
        RECT  0.22 0.84 0.52 1.12 ;
        RECT  0.22 0.96 0.84 1.12 ;
        RECT  0.54 0.96 0.70 2.26 ;
        RECT  0.54 1.98 0.90 2.26 ;
        RECT  2.04 0.84 2.32 1.12 ;
        RECT  1.78 0.96 2.32 1.12 ;
        RECT  1.66 1.98 1.94 2.26 ;
        RECT  1.78 0.96 1.94 2.64 ;
        RECT  1.78 2.48 2.60 2.64 ;
        RECT  2.32 2.48 2.60 2.76 ;
        RECT  2.90 0.68 3.18 0.96 ;
        RECT  2.90 0.80 3.45 0.96 ;
        RECT  3.29 1.12 4.25 1.28 ;
        RECT  4.09 1.12 4.25 1.78 ;
        RECT  4.09 1.50 4.37 1.78 ;
        RECT  3.29 0.80 3.45 2.26 ;
        RECT  3.28 1.98 3.56 2.26 ;
        RECT  5.13 0.96 5.54 1.24 ;
        RECT  5.38 1.45 5.82 1.73 ;
        RECT  5.38 0.96 5.54 1.82 ;
        RECT  4.53 1.66 5.56 1.82 ;
        RECT  5.40 1.45 5.56 2.24 ;
        RECT  4.53 1.66 4.69 2.24 ;
        RECT  4.36 1.96 4.69 2.24 ;
        RECT  5.40 1.96 5.68 2.24 ;
        RECT  5.88 0.74 6.16 1.24 ;
        RECT  5.98 1.46 6.90 1.62 ;
        RECT  6.62 1.40 6.90 1.68 ;
        RECT  5.98 0.74 6.14 2.46 ;
        RECT  5.88 1.96 6.16 2.46 ;
    END
END AND23OR3SP8V1_0

MACRO AND23OR3SP4V1_0
    CLASS CORE ;
    FOREIGN AND23OR3SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.40 1.14 1.82 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.40 0.38 1.82 ;
        END
    END IN1
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.40 1.62 1.82 ;
        END
    END IN3
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.10 1.40 2.38 1.82 ;
        END
    END IN4
    PIN IN5
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.85 1.40 3.13 1.82 ;
        END
    END IN5
    PIN IN6
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.61 1.52 3.93 1.82 ;
        RECT  3.61 1.46 3.89 1.82 ;
        END
    END IN6
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 13.33  LAYER ME1  ;
        ANTENNADIFFAREA 6.82  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.62  LAYER ME1  ;
        ANTENNAMAXAREACAR 21.52  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.96 1.96 7.48 2.12 ;
        RECT  7.32 1.08 7.48 2.12 ;
        RECT  6.96 1.08 7.48 1.24 ;
        RECT  6.96 1.96 7.24 2.46 ;
        RECT  6.96 0.74 7.24 1.24 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 7.60 3.48 ;
        RECT  7.14 2.88 7.42 3.48 ;
        RECT  6.44 1.96 6.72 2.46 ;
        RECT  6.50 1.96 6.66 3.48 ;
        RECT  4.88 2.24 5.16 2.52 ;
        RECT  4.95 2.24 5.11 3.48 ;
        RECT  3.84 2.24 4.12 2.52 ;
        RECT  3.90 2.24 4.06 3.48 ;
        RECT  2.76 1.98 3.04 2.26 ;
        RECT  2.82 1.98 2.98 3.48 ;
        RECT  1.14 1.98 1.42 2.26 ;
        RECT  1.20 1.98 1.36 3.48 ;
        RECT  0.10 1.98 0.38 2.26 ;
        RECT  0.16 1.98 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 7.60 0.28 ;
        RECT  7.14 -0.28 7.42 0.32 ;
        RECT  6.44 0.74 6.72 1.24 ;
        RECT  6.50 -0.28 6.66 1.24 ;
        RECT  3.85 0.68 4.13 0.96 ;
        RECT  3.91 -0.28 4.07 0.96 ;
        RECT  1.14 0.84 1.42 1.12 ;
        RECT  1.20 -0.28 1.36 1.12 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.44 0.38 0.72 ;
        RECT  0.22 0.44 0.38 1.12 ;
        RECT  0.22 0.84 0.52 1.12 ;
        RECT  0.22 0.96 0.84 1.12 ;
        RECT  0.54 0.96 0.70 2.26 ;
        RECT  0.54 1.98 0.90 2.26 ;
        RECT  2.04 0.84 2.32 1.12 ;
        RECT  1.78 0.96 2.32 1.12 ;
        RECT  1.66 1.98 1.94 2.26 ;
        RECT  1.78 0.96 1.94 2.64 ;
        RECT  1.78 2.48 2.60 2.64 ;
        RECT  2.32 2.48 2.60 2.76 ;
        RECT  2.90 0.68 3.18 0.96 ;
        RECT  2.90 0.80 3.45 0.96 ;
        RECT  3.29 1.12 4.25 1.28 ;
        RECT  4.09 1.12 4.25 1.78 ;
        RECT  4.09 1.50 4.37 1.78 ;
        RECT  3.29 0.80 3.45 2.26 ;
        RECT  3.28 1.98 3.56 2.26 ;
        RECT  5.13 0.96 5.54 1.24 ;
        RECT  5.38 1.45 5.82 1.73 ;
        RECT  5.38 0.96 5.54 1.82 ;
        RECT  4.53 1.66 5.56 1.82 ;
        RECT  5.40 1.45 5.56 2.24 ;
        RECT  4.53 1.66 4.69 2.24 ;
        RECT  4.36 1.96 4.69 2.24 ;
        RECT  5.40 1.96 5.68 2.24 ;
        RECT  5.88 0.84 6.16 1.24 ;
        RECT  5.98 1.46 6.90 1.62 ;
        RECT  6.62 1.40 6.90 1.68 ;
        RECT  5.98 0.84 6.14 2.36 ;
        RECT  5.88 1.96 6.16 2.36 ;
    END
END AND23OR3SP4V1_0

MACRO AND23OR3SP2V1_0
    CLASS CORE ;
    FOREIGN AND23OR3SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 10.05  LAYER ME1  ;
        ANTENNADIFFAREA 5.05  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.40  LAYER ME1  ;
        ANTENNAMAXAREACAR 24.92  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.40 1.96 5.68 2.24 ;
        RECT  5.40 1.66 5.56 2.24 ;
        RECT  5.32 0.96 5.48 1.82 ;
        RECT  4.53 1.66 5.56 1.82 ;
        RECT  5.13 0.96 5.48 1.24 ;
        RECT  4.36 1.96 4.69 2.24 ;
        RECT  4.53 1.66 4.69 2.24 ;
        END
    END OUT
    PIN IN6
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.61 1.52 3.93 1.82 ;
        RECT  3.61 1.46 3.89 1.82 ;
        END
    END IN6
    PIN IN5
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.85 1.40 3.13 1.82 ;
        END
    END IN5
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.10 1.40 2.38 1.82 ;
        END
    END IN4
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.40 1.62 1.82 ;
        END
    END IN3
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.40 0.38 1.82 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.40 1.14 1.82 ;
        END
    END IN2
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 6.00 0.28 ;
        RECT  5.54 -0.28 5.82 0.32 ;
        RECT  3.85 0.68 4.13 0.96 ;
        RECT  3.91 -0.28 4.07 0.96 ;
        RECT  1.14 0.84 1.42 1.12 ;
        RECT  1.20 -0.28 1.36 1.12 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 6.00 3.48 ;
        RECT  5.54 2.88 5.82 3.48 ;
        RECT  4.88 2.24 5.16 2.52 ;
        RECT  4.95 2.24 5.11 3.48 ;
        RECT  3.84 2.24 4.12 2.52 ;
        RECT  3.90 2.24 4.06 3.48 ;
        RECT  2.76 1.98 3.04 2.26 ;
        RECT  2.82 1.98 2.98 3.48 ;
        RECT  1.14 1.98 1.42 2.26 ;
        RECT  1.20 1.98 1.36 3.48 ;
        RECT  0.10 1.98 0.38 2.26 ;
        RECT  0.16 1.98 0.32 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.44 0.38 0.72 ;
        RECT  0.22 0.44 0.38 1.12 ;
        RECT  0.22 0.84 0.52 1.12 ;
        RECT  0.22 0.96 0.84 1.12 ;
        RECT  0.54 0.96 0.70 2.26 ;
        RECT  0.54 1.98 0.90 2.26 ;
        RECT  2.04 0.84 2.32 1.12 ;
        RECT  1.78 0.96 2.32 1.12 ;
        RECT  1.66 1.98 1.94 2.26 ;
        RECT  1.78 0.96 1.94 2.64 ;
        RECT  1.78 2.48 2.60 2.64 ;
        RECT  2.32 2.48 2.60 2.76 ;
        RECT  2.90 0.68 3.18 0.96 ;
        RECT  2.90 0.80 3.45 0.96 ;
        RECT  3.29 1.12 4.25 1.28 ;
        RECT  4.09 1.12 4.25 1.78 ;
        RECT  4.09 1.50 4.37 1.78 ;
        RECT  3.29 0.80 3.45 2.26 ;
        RECT  3.28 1.98 3.56 2.26 ;
    END
END AND23OR3SP2V1_0

MACRO AND23OR3SP1V1_0
    CLASS CORE ;
    FOREIGN AND23OR3SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 10.12  LAYER ME1  ;
        ANTENNADIFFAREA 4.27  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        ANTENNAMAXAREACAR 50.20  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.36 1.98 5.64 2.26 ;
        RECT  5.36 1.66 5.52 2.26 ;
        RECT  5.32 0.68 5.48 1.82 ;
        RECT  4.44 1.66 5.52 1.82 ;
        RECT  5.08 0.68 5.48 0.96 ;
        RECT  4.32 1.98 4.60 2.26 ;
        RECT  4.44 1.66 4.60 2.26 ;
        END
    END OUT
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.40 1.14 1.82 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.40 0.38 1.82 ;
        END
    END IN1
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.40 1.62 1.82 ;
        END
    END IN3
    PIN IN6
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.61 1.52 3.93 1.82 ;
        RECT  3.61 1.46 3.89 1.82 ;
        END
    END IN6
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.10 1.40 2.38 1.82 ;
        END
    END IN4
    PIN IN5
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.85 1.40 3.13 1.82 ;
        END
    END IN5
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 6.00 3.48 ;
        RECT  5.54 2.88 5.82 3.48 ;
        RECT  4.84 1.98 5.12 2.26 ;
        RECT  4.91 1.98 5.07 3.48 ;
        RECT  3.80 1.98 4.08 2.26 ;
        RECT  3.86 1.98 4.02 3.48 ;
        RECT  2.76 1.98 3.04 2.26 ;
        RECT  2.82 1.98 2.98 3.48 ;
        RECT  1.14 1.98 1.42 2.26 ;
        RECT  1.20 1.98 1.36 3.48 ;
        RECT  0.10 1.98 0.38 2.26 ;
        RECT  0.16 1.98 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 6.00 0.28 ;
        RECT  5.54 -0.28 5.82 0.32 ;
        RECT  3.80 0.68 4.08 0.96 ;
        RECT  3.86 -0.28 4.02 0.96 ;
        RECT  1.14 0.84 1.42 1.12 ;
        RECT  1.20 -0.28 1.36 1.12 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.44 0.38 0.72 ;
        RECT  0.22 0.44 0.38 1.12 ;
        RECT  0.22 0.84 0.52 1.12 ;
        RECT  0.22 0.96 0.84 1.12 ;
        RECT  0.54 0.96 0.70 2.26 ;
        RECT  0.54 1.98 0.90 2.26 ;
        RECT  2.04 0.84 2.32 1.12 ;
        RECT  1.78 0.96 2.32 1.12 ;
        RECT  1.66 1.98 1.94 2.26 ;
        RECT  1.78 0.96 1.94 2.64 ;
        RECT  1.78 2.48 2.60 2.64 ;
        RECT  2.32 2.48 2.60 2.76 ;
        RECT  2.90 0.68 3.18 0.96 ;
        RECT  2.90 0.80 3.45 0.96 ;
        RECT  3.29 1.12 4.32 1.28 ;
        RECT  4.04 1.12 4.32 1.40 ;
        RECT  3.29 0.80 3.45 2.26 ;
        RECT  3.28 1.98 3.56 2.26 ;
    END
END AND23OR3SP1V1_0

MACRO AND23NOR3SP8V1_0
    CLASS CORE ;
    FOREIGN AND23NOR3SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 14.72  LAYER ME1  ;
        ANTENNADIFFAREA 7.84  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.78  LAYER ME1  ;
        ANTENNAMAXAREACAR 18.93  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.42 1.98 7.70 2.26 ;
        RECT  6.38 1.08 7.70 1.24 ;
        RECT  7.42 0.64 7.70 1.24 ;
        RECT  6.38 1.98 7.70 2.14 ;
        RECT  6.38 1.98 6.68 2.26 ;
        RECT  6.52 0.64 6.68 2.26 ;
        RECT  6.38 0.64 6.68 1.24 ;
        END
    END OUT
    PIN IN6
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.66 1.40 3.94 1.82 ;
        END
    END IN6
    PIN IN5
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.86 1.40 3.14 1.82 ;
        END
    END IN5
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.40 1.62 1.82 ;
        END
    END IN3
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.10 1.40 2.38 1.82 ;
        END
    END IN4
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.40 0.38 1.82 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.40 1.14 1.82 ;
        END
    END IN2
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 8.40 3.48 ;
        RECT  7.94 2.88 8.22 3.48 ;
        RECT  7.94 2.30 8.22 2.58 ;
        RECT  8.00 2.30 8.16 3.48 ;
        RECT  6.90 2.30 7.18 2.58 ;
        RECT  6.96 2.30 7.12 3.48 ;
        RECT  5.86 2.30 6.14 2.58 ;
        RECT  5.92 2.30 6.08 3.48 ;
        RECT  4.78 1.98 5.06 2.26 ;
        RECT  4.84 1.98 5.00 3.48 ;
        RECT  3.78 1.98 4.06 2.26 ;
        RECT  3.84 1.98 4.00 3.48 ;
        RECT  2.84 2.10 3.00 3.48 ;
        RECT  2.50 2.10 3.00 2.26 ;
        RECT  2.50 1.98 2.78 2.26 ;
        RECT  1.14 1.98 1.42 2.26 ;
        RECT  1.20 1.98 1.36 3.48 ;
        RECT  0.10 1.98 0.38 2.26 ;
        RECT  0.16 1.98 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 8.40 0.28 ;
        RECT  7.94 0.64 8.22 1.24 ;
        RECT  7.94 -0.28 8.22 0.32 ;
        RECT  8.00 -0.28 8.16 1.24 ;
        RECT  6.90 0.64 7.18 0.92 ;
        RECT  6.96 -0.28 7.12 0.92 ;
        RECT  5.86 0.64 6.14 1.24 ;
        RECT  5.92 -0.28 6.08 1.24 ;
        RECT  2.74 0.96 3.02 1.24 ;
        RECT  2.80 -0.28 2.96 1.24 ;
        RECT  1.08 0.84 1.36 1.12 ;
        RECT  1.14 -0.28 1.30 1.12 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.44 0.38 0.72 ;
        RECT  0.22 0.44 0.38 1.12 ;
        RECT  0.22 0.84 0.52 1.12 ;
        RECT  0.22 0.96 0.70 1.12 ;
        RECT  0.54 0.96 0.70 2.26 ;
        RECT  0.54 1.98 0.90 2.26 ;
        RECT  2.12 0.84 2.40 1.12 ;
        RECT  1.78 0.96 2.40 1.12 ;
        RECT  1.66 1.98 1.94 2.26 ;
        RECT  1.78 0.96 1.94 2.64 ;
        RECT  1.78 2.48 2.68 2.64 ;
        RECT  2.40 2.48 2.68 2.76 ;
        RECT  3.78 0.58 4.06 0.86 ;
        RECT  3.64 0.96 3.94 1.24 ;
        RECT  3.78 0.58 3.94 1.24 ;
        RECT  3.34 1.08 3.94 1.24 ;
        RECT  3.34 1.08 3.50 2.26 ;
        RECT  3.26 1.98 3.54 2.26 ;
        RECT  4.54 0.96 4.82 1.24 ;
        RECT  4.60 0.96 4.76 1.82 ;
        RECT  6.08 1.54 6.36 1.82 ;
        RECT  4.38 1.66 6.36 1.82 ;
        RECT  5.30 1.66 5.46 2.26 ;
        RECT  4.38 1.66 4.54 2.26 ;
        RECT  4.26 1.98 4.54 2.26 ;
        RECT  5.30 1.98 5.58 2.26 ;
    END
END AND23NOR3SP8V1_0

MACRO AND23NOR3SP4V1_0
    CLASS CORE ;
    FOREIGN AND23NOR3SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.40 1.14 1.82 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.40 0.38 1.82 ;
        END
    END IN1
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.10 1.40 2.38 1.82 ;
        END
    END IN4
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.40 1.62 1.82 ;
        END
    END IN3
    PIN IN5
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.86 1.40 3.14 1.82 ;
        END
    END IN5
    PIN IN6
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.66 1.40 3.94 1.82 ;
        END
    END IN6
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 12.70  LAYER ME1  ;
        ANTENNADIFFAREA 6.62  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER ME1  ;
        ANTENNAMAXAREACAR 25.94  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.38 1.98 6.68 2.26 ;
        RECT  6.52 0.64 6.68 2.26 ;
        RECT  6.38 0.64 6.68 1.24 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 7.60 3.48 ;
        RECT  6.98 2.88 7.42 3.48 ;
        RECT  6.90 2.30 7.18 2.58 ;
        RECT  6.98 2.30 7.14 3.48 ;
        RECT  5.86 2.30 6.14 2.58 ;
        RECT  5.92 2.30 6.08 3.48 ;
        RECT  4.78 1.98 5.06 2.26 ;
        RECT  4.84 1.98 5.00 3.48 ;
        RECT  3.78 1.98 4.06 2.26 ;
        RECT  3.84 1.98 4.00 3.48 ;
        RECT  2.84 2.10 3.00 3.48 ;
        RECT  2.50 2.10 3.00 2.26 ;
        RECT  2.50 1.98 2.78 2.26 ;
        RECT  1.14 1.98 1.42 2.26 ;
        RECT  1.20 1.98 1.36 3.48 ;
        RECT  0.10 1.98 0.38 2.26 ;
        RECT  0.16 1.98 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 7.60 0.28 ;
        RECT  6.98 -0.28 7.42 0.32 ;
        RECT  6.90 0.64 7.18 1.24 ;
        RECT  6.98 -0.28 7.14 1.24 ;
        RECT  5.86 0.64 6.14 1.24 ;
        RECT  5.92 -0.28 6.08 1.24 ;
        RECT  2.74 0.96 3.02 1.24 ;
        RECT  2.80 -0.28 2.96 1.24 ;
        RECT  1.08 0.84 1.36 1.12 ;
        RECT  1.14 -0.28 1.30 1.12 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.44 0.38 0.72 ;
        RECT  0.22 0.44 0.38 1.12 ;
        RECT  0.22 0.84 0.52 1.12 ;
        RECT  0.22 0.96 0.70 1.12 ;
        RECT  0.54 0.96 0.70 2.26 ;
        RECT  0.54 1.98 0.90 2.26 ;
        RECT  2.12 0.84 2.40 1.12 ;
        RECT  1.78 0.96 2.40 1.12 ;
        RECT  1.66 1.98 1.94 2.26 ;
        RECT  1.78 0.96 1.94 2.64 ;
        RECT  1.78 2.48 2.68 2.64 ;
        RECT  2.40 2.48 2.68 2.76 ;
        RECT  3.78 0.58 4.06 0.86 ;
        RECT  3.64 0.96 3.94 1.24 ;
        RECT  3.78 0.58 3.94 1.24 ;
        RECT  3.34 1.08 3.94 1.24 ;
        RECT  3.34 1.08 3.50 2.26 ;
        RECT  3.26 1.98 3.54 2.26 ;
        RECT  4.54 0.96 4.82 1.24 ;
        RECT  4.60 0.96 4.76 1.82 ;
        RECT  6.08 1.54 6.36 1.82 ;
        RECT  4.38 1.66 6.36 1.82 ;
        RECT  5.30 1.66 5.46 2.26 ;
        RECT  4.38 1.66 4.54 2.26 ;
        RECT  4.26 1.98 4.54 2.26 ;
        RECT  5.30 1.98 5.58 2.26 ;
    END
END AND23NOR3SP4V1_0

MACRO AND23NOR3SP2V1_0
    CLASS CORE ;
    FOREIGN AND23NOR3SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 11.44  LAYER ME1  ;
        ANTENNADIFFAREA 5.50  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.35  LAYER ME1  ;
        ANTENNAMAXAREACAR 33.12  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.38 1.98 6.68 2.26 ;
        RECT  6.52 0.64 6.68 2.26 ;
        RECT  6.38 0.64 6.68 1.24 ;
        END
    END OUT
    PIN IN6
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.66 1.40 3.94 1.82 ;
        END
    END IN6
    PIN IN5
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.86 1.40 3.14 1.82 ;
        END
    END IN5
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.40 1.62 1.82 ;
        END
    END IN3
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.10 1.40 2.38 1.82 ;
        END
    END IN4
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.40 0.38 1.82 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.40 1.14 1.82 ;
        END
    END IN2
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 6.80 0.28 ;
        RECT  6.34 -0.28 6.62 0.32 ;
        RECT  5.86 0.64 6.14 1.24 ;
        RECT  5.92 -0.28 6.08 1.24 ;
        RECT  2.74 0.96 3.02 1.24 ;
        RECT  2.80 -0.28 2.96 1.24 ;
        RECT  1.08 0.84 1.36 1.12 ;
        RECT  1.14 -0.28 1.30 1.12 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 6.80 3.48 ;
        RECT  6.34 2.88 6.62 3.48 ;
        RECT  5.86 2.30 6.14 2.58 ;
        RECT  5.92 2.30 6.08 3.48 ;
        RECT  4.78 1.98 5.06 2.26 ;
        RECT  4.84 1.98 5.00 3.48 ;
        RECT  3.78 1.98 4.06 2.26 ;
        RECT  3.84 1.98 4.00 3.48 ;
        RECT  2.84 2.10 3.00 3.48 ;
        RECT  2.50 2.10 3.00 2.26 ;
        RECT  2.50 1.98 2.78 2.26 ;
        RECT  1.14 1.98 1.42 2.26 ;
        RECT  1.20 1.98 1.36 3.48 ;
        RECT  0.10 1.98 0.38 2.26 ;
        RECT  0.16 1.98 0.32 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.44 0.38 0.72 ;
        RECT  0.22 0.44 0.38 1.12 ;
        RECT  0.22 0.84 0.52 1.12 ;
        RECT  0.22 0.96 0.70 1.12 ;
        RECT  0.54 0.96 0.70 2.26 ;
        RECT  0.54 1.98 0.90 2.26 ;
        RECT  2.12 0.84 2.40 1.12 ;
        RECT  1.78 0.96 2.40 1.12 ;
        RECT  1.66 1.98 1.94 2.26 ;
        RECT  1.78 0.96 1.94 2.64 ;
        RECT  1.78 2.48 2.68 2.64 ;
        RECT  2.40 2.48 2.68 2.76 ;
        RECT  3.78 0.58 4.06 0.86 ;
        RECT  3.64 0.96 3.94 1.24 ;
        RECT  3.78 0.58 3.94 1.24 ;
        RECT  3.34 1.08 3.94 1.24 ;
        RECT  3.34 1.08 3.50 2.26 ;
        RECT  3.26 1.98 3.54 2.26 ;
        RECT  4.54 0.96 4.82 1.24 ;
        RECT  4.60 0.96 4.76 1.82 ;
        RECT  6.08 1.54 6.36 1.82 ;
        RECT  4.38 1.66 6.36 1.82 ;
        RECT  5.30 1.66 5.46 2.26 ;
        RECT  4.38 1.66 4.54 2.26 ;
        RECT  4.26 1.98 4.54 2.26 ;
        RECT  5.30 1.98 5.58 2.26 ;
    END
END AND23NOR3SP2V1_0

MACRO AND23NOR3SP1V1_0
    CLASS CORE ;
    FOREIGN AND23NOR3SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 11.46  LAYER ME1  ;
        ANTENNADIFFAREA 5.04  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.27  LAYER ME1  ;
        ANTENNAMAXAREACAR 42.63  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.34 1.98 6.68 2.26 ;
        RECT  6.52 0.96 6.68 2.26 ;
        RECT  6.34 0.96 6.68 1.24 ;
        END
    END OUT
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.40 1.14 1.82 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.40 0.38 1.82 ;
        END
    END IN1
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.10 1.40 2.38 1.82 ;
        END
    END IN4
    PIN IN5
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.86 1.40 3.14 1.82 ;
        END
    END IN5
    PIN IN6
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.66 1.40 3.94 1.82 ;
        END
    END IN6
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.40 1.62 1.82 ;
        END
    END IN3
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 6.80 3.48 ;
        RECT  6.34 2.88 6.62 3.48 ;
        RECT  5.82 1.98 6.10 2.26 ;
        RECT  5.88 1.98 6.04 3.48 ;
        RECT  4.78 1.98 5.06 2.26 ;
        RECT  4.84 1.98 5.00 3.48 ;
        RECT  3.78 1.98 4.06 2.26 ;
        RECT  3.84 1.98 4.00 3.48 ;
        RECT  2.84 2.10 3.00 3.48 ;
        RECT  2.50 2.10 3.00 2.26 ;
        RECT  2.50 1.98 2.78 2.26 ;
        RECT  1.14 1.98 1.42 2.26 ;
        RECT  1.20 1.98 1.36 3.48 ;
        RECT  0.10 1.98 0.38 2.26 ;
        RECT  0.17 1.98 0.33 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 6.80 0.28 ;
        RECT  6.34 -0.28 6.62 0.32 ;
        RECT  5.82 0.96 6.10 1.24 ;
        RECT  5.88 -0.28 6.04 1.24 ;
        RECT  2.74 0.96 3.02 1.24 ;
        RECT  2.80 -0.28 2.96 1.24 ;
        RECT  1.08 0.84 1.36 1.12 ;
        RECT  1.14 -0.28 1.30 1.12 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.44 0.38 0.72 ;
        RECT  0.22 0.44 0.38 1.12 ;
        RECT  0.22 0.84 0.52 1.12 ;
        RECT  0.22 0.96 0.70 1.12 ;
        RECT  0.54 0.96 0.70 2.26 ;
        RECT  0.54 1.98 0.90 2.26 ;
        RECT  2.12 0.84 2.40 1.12 ;
        RECT  1.78 0.96 2.40 1.12 ;
        RECT  1.66 1.98 1.94 2.26 ;
        RECT  1.78 0.96 1.94 2.64 ;
        RECT  1.78 2.48 2.68 2.64 ;
        RECT  2.40 2.48 2.68 2.76 ;
        RECT  3.78 0.58 4.06 0.86 ;
        RECT  3.64 0.96 3.94 1.24 ;
        RECT  3.78 0.58 3.94 1.24 ;
        RECT  3.34 1.08 3.94 1.24 ;
        RECT  3.34 1.08 3.50 2.26 ;
        RECT  3.26 1.98 3.54 2.26 ;
        RECT  4.54 0.96 4.82 1.24 ;
        RECT  4.60 0.96 4.76 1.82 ;
        RECT  6.08 1.54 6.36 1.82 ;
        RECT  4.38 1.66 6.36 1.82 ;
        RECT  5.30 1.66 5.46 2.26 ;
        RECT  4.38 1.66 4.54 2.26 ;
        RECT  4.26 1.98 4.54 2.26 ;
        RECT  5.30 1.98 5.58 2.26 ;
    END
END AND23NOR3SP1V1_0

MACRO AND22OR2SP8V1_0
    CLASS CORE ;
    FOREIGN AND22OR2SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.66 1.40 1.96 1.75 ;
        END
    END IN3
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.12 1.40 2.45 1.74 ;
        END
    END IN4
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 14.42  LAYER ME1  ;
        ANTENNADIFFAREA 7.87  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER ME1  ;
        ANTENNAMAXAREACAR 12.52  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.52 2.23 6.80 2.51 ;
        RECT  6.52 0.96 6.80 1.24 ;
        RECT  6.52 2.06 6.68 2.51 ;
        RECT  5.54 1.52 6.68 1.68 ;
        RECT  6.52 0.96 6.68 1.68 ;
        RECT  3.52 2.06 6.68 2.22 ;
        RECT  5.48 2.06 5.76 2.51 ;
        RECT  5.48 0.96 5.76 1.24 ;
        RECT  5.54 0.96 5.70 2.51 ;
        RECT  4.44 2.06 4.72 2.51 ;
        RECT  3.40 2.23 3.68 2.51 ;
        RECT  3.52 2.06 3.68 2.51 ;
        END
    END OUT
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.90 1.32 1.18 1.74 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.46 0.93 0.74 1.35 ;
        END
    END IN1
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 7.60 0.28 ;
        RECT  7.14 -0.28 7.42 0.32 ;
        RECT  4.44 0.64 4.72 0.92 ;
        RECT  4.49 -0.28 4.65 0.92 ;
        RECT  3.40 0.64 3.68 0.92 ;
        RECT  3.46 -0.28 3.62 0.92 ;
        RECT  2.40 0.96 2.68 1.24 ;
        RECT  2.46 -0.28 2.62 1.24 ;
        RECT  1.16 0.49 1.44 0.77 ;
        RECT  1.22 -0.28 1.38 0.77 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 7.60 3.48 ;
        RECT  7.10 2.88 7.42 3.48 ;
        RECT  7.04 2.38 7.32 2.66 ;
        RECT  7.10 2.38 7.26 3.48 ;
        RECT  6.00 2.38 6.28 2.66 ;
        RECT  6.06 2.38 6.22 3.48 ;
        RECT  4.96 2.38 5.24 2.66 ;
        RECT  5.02 2.38 5.18 3.48 ;
        RECT  3.92 2.38 4.20 2.66 ;
        RECT  3.98 2.38 4.14 3.48 ;
        RECT  2.88 2.38 3.16 2.66 ;
        RECT  2.94 2.38 3.10 3.48 ;
        RECT  2.40 2.23 2.68 2.51 ;
        RECT  2.46 2.23 2.62 3.48 ;
        RECT  1.36 2.23 1.64 2.51 ;
        RECT  1.42 2.23 1.58 3.48 ;
        RECT  0.32 2.23 0.60 2.51 ;
        RECT  0.38 2.23 0.54 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.14 0.49 0.60 0.77 ;
        RECT  0.14 0.49 0.30 1.77 ;
        RECT  0.10 1.49 0.38 1.77 ;
        RECT  0.22 1.49 0.38 2.07 ;
        RECT  0.22 1.91 1.00 2.07 ;
        RECT  0.84 1.91 1.00 2.51 ;
        RECT  0.84 2.23 1.12 2.51 ;
        RECT  1.34 0.96 1.79 1.24 ;
        RECT  5.10 1.46 5.38 1.74 ;
        RECT  2.76 1.58 5.38 1.74 ;
        RECT  1.34 0.96 1.50 2.07 ;
        RECT  2.76 1.58 2.92 2.07 ;
        RECT  1.34 1.91 2.92 2.07 ;
        RECT  1.88 1.91 2.04 2.51 ;
        RECT  1.88 2.23 2.16 2.51 ;
        RECT  4.96 0.64 7.32 0.80 ;
        RECT  2.88 0.64 3.16 1.24 ;
        RECT  3.92 0.64 4.20 1.24 ;
        RECT  4.96 0.64 5.24 1.24 ;
        RECT  2.88 1.08 5.24 1.24 ;
        RECT  6.00 0.64 6.28 1.24 ;
        RECT  7.04 0.64 7.32 1.24 ;
    END
END AND22OR2SP8V1_0

MACRO AND22OR2SP4V1_0
    CLASS CORE ;
    FOREIGN AND22OR2SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.60 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.46 0.93 0.74 1.35 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.90 1.32 1.18 1.74 ;
        END
    END IN2
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 9.74  LAYER ME1  ;
        ANTENNADIFFAREA 5.31  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.58  LAYER ME1  ;
        ANTENNAMAXAREACAR 16.92  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.44 2.06 4.72 2.51 ;
        RECT  4.56 0.96 4.72 2.51 ;
        RECT  4.44 0.96 4.72 1.24 ;
        RECT  3.52 2.06 4.72 2.22 ;
        RECT  3.40 2.23 3.68 2.51 ;
        RECT  3.52 2.06 3.68 2.51 ;
        END
    END OUT
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.12 1.40 2.45 1.74 ;
        END
    END IN4
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.66 1.40 1.96 1.75 ;
        END
    END IN3
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 5.60 3.48 ;
        RECT  5.02 2.88 5.42 3.48 ;
        RECT  4.96 2.38 5.24 2.66 ;
        RECT  5.02 2.38 5.18 3.48 ;
        RECT  3.92 2.38 4.20 2.66 ;
        RECT  3.98 2.38 4.14 3.48 ;
        RECT  2.88 2.38 3.16 2.66 ;
        RECT  2.94 2.38 3.10 3.48 ;
        RECT  2.40 2.23 2.68 2.51 ;
        RECT  2.46 2.23 2.62 3.48 ;
        RECT  1.36 2.23 1.64 2.51 ;
        RECT  1.42 2.23 1.58 3.48 ;
        RECT  0.32 2.23 0.60 2.51 ;
        RECT  0.38 2.23 0.54 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 5.60 0.28 ;
        RECT  5.14 -0.28 5.42 0.32 ;
        RECT  3.40 0.64 3.68 0.92 ;
        RECT  3.46 -0.28 3.62 0.92 ;
        RECT  2.40 0.96 2.68 1.24 ;
        RECT  2.46 -0.28 2.62 1.24 ;
        RECT  1.16 0.49 1.44 0.77 ;
        RECT  1.22 -0.28 1.38 0.77 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.14 0.49 0.60 0.77 ;
        RECT  0.14 0.49 0.30 1.77 ;
        RECT  0.10 1.49 0.38 1.77 ;
        RECT  0.22 1.49 0.38 2.07 ;
        RECT  0.22 1.91 1.00 2.07 ;
        RECT  0.84 1.91 1.00 2.51 ;
        RECT  0.84 2.23 1.12 2.51 ;
        RECT  1.34 0.96 1.79 1.24 ;
        RECT  4.06 1.46 4.34 1.74 ;
        RECT  2.76 1.58 4.34 1.74 ;
        RECT  1.34 0.96 1.50 2.07 ;
        RECT  2.76 1.58 2.92 2.07 ;
        RECT  1.34 1.91 2.92 2.07 ;
        RECT  1.88 1.91 2.04 2.51 ;
        RECT  1.88 2.23 2.16 2.51 ;
        RECT  3.92 0.64 5.24 0.80 ;
        RECT  2.88 0.64 3.16 1.24 ;
        RECT  3.92 0.64 4.20 1.24 ;
        RECT  2.88 1.08 4.20 1.24 ;
        RECT  4.96 0.64 5.24 1.24 ;
    END
END AND22OR2SP4V1_0

MACRO AND22OR2SP2V1_0
    CLASS CORE ;
    FOREIGN AND22OR2SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.66 1.40 1.96 1.75 ;
        END
    END IN3
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.12 1.40 2.45 1.74 ;
        END
    END IN4
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 7.39  LAYER ME1  ;
        ANTENNADIFFAREA 3.58  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.29  LAYER ME1  ;
        ANTENNAMAXAREACAR 25.66  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.12 1.91 3.88 2.07 ;
        RECT  3.72 0.64 3.88 2.07 ;
        RECT  3.28 0.64 3.88 1.24 ;
        RECT  2.96 2.23 3.28 2.51 ;
        RECT  3.12 1.91 3.28 2.51 ;
        END
    END OUT
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.90 1.32 1.18 1.74 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.46 0.93 0.74 1.35 ;
        END
    END IN1
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.00 0.28 ;
        RECT  3.54 -0.28 3.82 0.32 ;
        RECT  2.44 0.64 2.72 1.24 ;
        RECT  2.50 -0.28 2.66 1.24 ;
        RECT  1.16 0.49 1.44 0.77 ;
        RECT  1.22 -0.28 1.38 0.77 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.00 3.48 ;
        RECT  3.54 2.88 3.82 3.48 ;
        RECT  3.48 2.38 3.76 2.66 ;
        RECT  3.54 2.38 3.70 3.48 ;
        RECT  2.44 2.38 2.72 2.66 ;
        RECT  2.50 2.38 2.66 3.48 ;
        RECT  1.36 2.23 1.64 2.51 ;
        RECT  1.42 2.23 1.58 3.48 ;
        RECT  0.32 2.23 0.60 2.51 ;
        RECT  0.38 2.23 0.54 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.14 0.49 0.60 0.77 ;
        RECT  0.14 0.49 0.30 1.77 ;
        RECT  0.10 1.49 0.38 1.77 ;
        RECT  0.22 1.49 0.38 2.07 ;
        RECT  0.22 1.91 1.00 2.07 ;
        RECT  0.84 1.91 1.00 2.51 ;
        RECT  0.84 2.23 1.12 2.51 ;
        RECT  1.34 0.96 1.79 1.24 ;
        RECT  3.10 1.46 3.38 1.74 ;
        RECT  2.80 1.58 3.38 1.74 ;
        RECT  1.34 0.96 1.50 2.07 ;
        RECT  2.80 1.58 2.96 2.07 ;
        RECT  1.34 1.91 2.96 2.07 ;
        RECT  1.88 1.91 2.04 2.51 ;
        RECT  1.88 2.23 2.16 2.51 ;
    END
END AND22OR2SP2V1_0

MACRO AND22OR2SP1V1_0
    CLASS CORE ;
    FOREIGN AND22OR2SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.00 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 6.69  LAYER ME1  ;
        ANTENNADIFFAREA 2.93  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.13  LAYER ME1  ;
        ANTENNAMAXAREACAR 49.78  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.12 1.91 3.88 2.07 ;
        RECT  3.72 0.96 3.88 2.07 ;
        RECT  3.24 0.96 3.88 1.24 ;
        RECT  2.92 2.23 3.28 2.51 ;
        RECT  3.12 1.91 3.28 2.51 ;
        END
    END OUT
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.90 1.32 1.18 1.74 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.46 0.93 0.74 1.35 ;
        END
    END IN1
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.66 1.40 1.96 1.75 ;
        END
    END IN3
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.12 1.40 2.45 1.74 ;
        END
    END IN4
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.00 0.28 ;
        RECT  3.54 -0.28 3.82 0.32 ;
        RECT  2.40 0.96 2.68 1.24 ;
        RECT  2.46 -0.28 2.62 1.24 ;
        RECT  1.16 0.49 1.44 0.77 ;
        RECT  1.22 -0.28 1.38 0.77 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.00 3.48 ;
        RECT  3.50 2.88 3.82 3.48 ;
        RECT  3.44 2.23 3.72 2.51 ;
        RECT  3.50 2.23 3.66 3.48 ;
        RECT  2.40 2.23 2.68 2.51 ;
        RECT  2.46 2.23 2.62 3.48 ;
        RECT  1.36 2.23 1.64 2.51 ;
        RECT  1.42 2.23 1.58 3.48 ;
        RECT  0.32 2.23 0.60 2.51 ;
        RECT  0.38 2.23 0.54 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.14 0.49 0.60 0.77 ;
        RECT  0.14 0.49 0.30 1.77 ;
        RECT  0.10 1.49 0.38 1.77 ;
        RECT  0.22 1.49 0.38 2.07 ;
        RECT  0.22 1.91 1.00 2.07 ;
        RECT  0.84 1.91 1.00 2.51 ;
        RECT  0.84 2.23 1.12 2.51 ;
        RECT  1.34 0.96 1.79 1.24 ;
        RECT  3.06 1.46 3.34 1.74 ;
        RECT  2.80 1.58 3.34 1.74 ;
        RECT  1.34 0.96 1.50 2.07 ;
        RECT  2.80 1.58 2.96 2.07 ;
        RECT  1.34 1.91 2.96 2.07 ;
        RECT  1.88 1.91 2.04 2.51 ;
        RECT  1.88 2.23 2.16 2.51 ;
    END
END AND22OR2SP1V1_0

MACRO AND22NOR2SP8V1_0
    CLASS CORE ;
    FOREIGN AND22NOR2SP8V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 12.10  LAYER ME1  ;
        ANTENNADIFFAREA 6.07  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.71  LAYER ME1  ;
        ANTENNAMAXAREACAR 17.03  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.30 1.97 5.58 2.57 ;
        RECT  5.30 0.64 5.58 1.24 ;
        RECT  5.30 0.64 5.46 2.57 ;
        RECT  4.46 1.52 5.46 1.68 ;
        RECT  4.26 1.97 4.62 2.57 ;
        RECT  4.46 0.64 4.62 2.57 ;
        RECT  4.26 0.64 4.62 1.24 ;
        END
    END OUT
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.10 1.40 2.38 1.82 ;
        END
    END IN4
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.40 1.62 1.82 ;
        END
    END IN3
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.40 0.38 1.82 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.46 1.14 1.86 ;
        END
    END IN2
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 6.40 0.28 ;
        RECT  5.88 -0.28 6.22 0.32 ;
        RECT  5.82 0.64 6.10 1.24 ;
        RECT  5.88 -0.28 6.04 1.24 ;
        RECT  4.78 0.64 5.06 1.24 ;
        RECT  4.84 -0.28 5.00 1.24 ;
        RECT  3.74 0.64 4.02 1.24 ;
        RECT  3.80 -0.28 3.96 1.24 ;
        RECT  1.16 0.96 1.44 1.24 ;
        RECT  1.22 -0.28 1.38 1.24 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 6.40 3.48 ;
        RECT  5.88 2.88 6.22 3.48 ;
        RECT  5.82 1.97 6.10 2.57 ;
        RECT  5.88 1.97 6.04 3.48 ;
        RECT  4.78 1.97 5.06 2.57 ;
        RECT  4.84 1.97 5.00 3.48 ;
        RECT  3.74 1.97 4.02 2.57 ;
        RECT  3.80 1.97 3.96 3.48 ;
        RECT  2.66 1.97 2.94 2.25 ;
        RECT  2.72 1.97 2.88 3.48 ;
        RECT  2.18 2.02 2.46 2.30 ;
        RECT  2.24 2.02 2.40 3.48 ;
        RECT  1.14 2.02 1.42 2.30 ;
        RECT  1.20 2.02 1.36 3.48 ;
        RECT  0.10 2.02 0.38 2.30 ;
        RECT  0.16 2.02 0.32 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.44 0.38 0.72 ;
        RECT  0.22 0.44 0.38 1.24 ;
        RECT  0.22 0.96 0.52 1.24 ;
        RECT  0.22 1.08 0.70 1.24 ;
        RECT  0.54 1.08 0.70 2.30 ;
        RECT  0.54 2.02 0.90 2.30 ;
        RECT  2.08 0.96 2.36 1.24 ;
        RECT  1.78 1.08 2.70 1.24 ;
        RECT  2.54 1.08 2.70 1.74 ;
        RECT  2.54 1.46 2.94 1.74 ;
        RECT  1.78 1.08 1.94 2.30 ;
        RECT  1.66 2.02 1.94 2.30 ;
        RECT  2.86 0.68 3.26 0.96 ;
        RECT  3.10 1.52 4.25 1.68 ;
        RECT  3.97 1.46 4.25 1.74 ;
        RECT  3.10 0.68 3.26 2.25 ;
        RECT  3.10 1.97 3.46 2.25 ;
    END
END AND22NOR2SP8V1_0

MACRO AND22NOR2SP4V1_0
    CLASS CORE ;
    FOREIGN AND22NOR2SP4V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.20 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.46 1.14 1.86 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.40 0.38 1.82 ;
        END
    END IN1
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.40 1.62 1.82 ;
        END
    END IN3
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.10 1.40 2.38 1.82 ;
        END
    END IN4
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 9.75  LAYER ME1  ;
        ANTENNADIFFAREA 4.73  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.42  LAYER ME1  ;
        ANTENNAMAXAREACAR 23.08  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.46 1.52 4.68 1.68 ;
        RECT  4.26 1.97 4.62 2.57 ;
        RECT  4.46 0.64 4.62 2.57 ;
        RECT  4.26 0.64 4.62 1.24 ;
        END
    END OUT
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 5.20 3.48 ;
        RECT  4.78 1.97 5.06 2.57 ;
        RECT  4.74 2.88 5.02 3.48 ;
        RECT  4.84 1.97 5.00 3.48 ;
        RECT  3.74 1.97 4.02 2.57 ;
        RECT  3.80 1.97 3.96 3.48 ;
        RECT  2.66 1.97 2.94 2.25 ;
        RECT  2.72 1.97 2.88 3.48 ;
        RECT  2.18 2.02 2.46 2.30 ;
        RECT  2.24 2.02 2.40 3.48 ;
        RECT  1.14 2.02 1.42 2.30 ;
        RECT  1.20 2.02 1.36 3.48 ;
        RECT  0.10 2.02 0.38 2.30 ;
        RECT  0.16 2.02 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 5.20 0.28 ;
        RECT  4.78 0.64 5.06 1.24 ;
        RECT  4.74 -0.28 5.02 0.32 ;
        RECT  4.84 -0.28 5.00 1.24 ;
        RECT  3.74 0.64 4.02 1.24 ;
        RECT  3.80 -0.28 3.96 1.24 ;
        RECT  1.16 0.96 1.44 1.24 ;
        RECT  1.22 -0.28 1.38 1.24 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.44 0.38 0.72 ;
        RECT  0.22 0.44 0.38 1.24 ;
        RECT  0.22 0.96 0.52 1.24 ;
        RECT  0.22 1.08 0.70 1.24 ;
        RECT  0.54 1.08 0.70 2.30 ;
        RECT  0.54 2.02 0.90 2.30 ;
        RECT  2.08 0.96 2.36 1.24 ;
        RECT  1.78 1.08 2.70 1.24 ;
        RECT  2.54 1.08 2.70 1.74 ;
        RECT  2.54 1.46 2.94 1.74 ;
        RECT  1.78 1.08 1.94 2.30 ;
        RECT  1.66 2.02 1.94 2.30 ;
        RECT  2.86 0.68 3.26 0.96 ;
        RECT  3.10 1.52 4.25 1.68 ;
        RECT  3.97 1.46 4.25 1.74 ;
        RECT  3.10 0.68 3.26 2.25 ;
        RECT  3.10 1.97 3.46 2.25 ;
    END
END AND22NOR2SP4V1_0

MACRO AND22NOR2SP2V1_0
    CLASS CORE ;
    FOREIGN AND22NOR2SP2V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 8.93  LAYER ME1  ;
        ANTENNADIFFAREA 3.89  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.28  LAYER ME1  ;
        ANTENNAMAXAREACAR 32.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.26 1.97 4.68 2.57 ;
        RECT  4.52 0.64 4.68 2.57 ;
        RECT  4.26 0.64 4.68 1.24 ;
        END
    END OUT
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.10 1.40 2.38 1.82 ;
        END
    END IN4
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.40 1.62 1.82 ;
        END
    END IN3
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.10 1.40 0.38 1.82 ;
        END
    END IN1
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.46 1.14 1.86 ;
        END
    END IN2
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.80 0.28 ;
        RECT  4.34 -0.28 4.62 0.32 ;
        RECT  3.74 0.64 4.02 1.24 ;
        RECT  3.80 -0.28 3.96 1.24 ;
        RECT  1.16 0.96 1.44 1.24 ;
        RECT  1.22 -0.28 1.38 1.24 ;
        END
    END GND!
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.80 3.48 ;
        RECT  4.34 2.88 4.62 3.48 ;
        RECT  3.74 1.97 4.02 2.57 ;
        RECT  3.80 1.97 3.96 3.48 ;
        RECT  2.66 1.97 2.94 2.25 ;
        RECT  2.72 1.97 2.88 3.48 ;
        RECT  2.18 2.02 2.46 2.30 ;
        RECT  2.24 2.02 2.40 3.48 ;
        RECT  1.14 2.02 1.42 2.30 ;
        RECT  1.20 2.02 1.36 3.48 ;
        RECT  0.10 2.02 0.38 2.30 ;
        RECT  0.16 2.02 0.32 3.48 ;
        END
    END VDD!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.44 0.38 0.72 ;
        RECT  0.22 0.44 0.38 1.24 ;
        RECT  0.22 0.96 0.52 1.24 ;
        RECT  0.22 1.08 0.70 1.24 ;
        RECT  0.54 1.08 0.70 2.30 ;
        RECT  0.54 2.02 0.90 2.30 ;
        RECT  2.08 0.96 2.36 1.24 ;
        RECT  1.78 1.08 2.70 1.24 ;
        RECT  2.54 1.08 2.70 1.74 ;
        RECT  2.54 1.46 2.94 1.74 ;
        RECT  1.78 1.08 1.94 2.30 ;
        RECT  1.66 2.02 1.94 2.30 ;
        RECT  2.86 0.68 3.26 0.96 ;
        RECT  3.10 1.52 4.25 1.68 ;
        RECT  3.97 1.46 4.25 1.74 ;
        RECT  3.10 0.68 3.26 2.25 ;
        RECT  3.10 1.97 3.46 2.25 ;
    END
END AND22NOR2SP2V1_0

MACRO AND22NOR2SP1V1_0
    CLASS CORE ;
    FOREIGN AND22NOR2SP1V1_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.80 BY 3.20 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN OUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALAREA 8.18  LAYER ME1  ;
        ANTENNADIFFAREA 3.43  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.20  LAYER ME1  ;
        ANTENNAMAXAREACAR 40.60  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.22 1.97 4.68 2.13 ;
        RECT  4.52 0.80 4.68 2.13 ;
        RECT  4.22 0.80 4.68 0.96 ;
        RECT  4.22 1.97 4.50 2.25 ;
        RECT  4.22 0.68 4.50 0.96 ;
        END
    END OUT
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.86 1.46 1.14 1.86 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.08 1.40 0.38 1.82 ;
        END
    END IN1
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.10 1.40 2.38 1.82 ;
        END
    END IN4
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.07  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.30 1.40 1.62 1.82 ;
        END
    END IN3
    PIN VDD!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 2.92 4.80 3.48 ;
        RECT  4.34 2.88 4.62 3.48 ;
        RECT  3.70 1.97 3.98 2.25 ;
        RECT  3.76 1.97 3.92 3.48 ;
        RECT  2.66 1.97 2.94 2.25 ;
        RECT  2.72 1.97 2.88 3.48 ;
        RECT  2.18 2.02 2.46 2.30 ;
        RECT  2.24 2.02 2.40 3.48 ;
        RECT  1.14 2.02 1.42 2.30 ;
        RECT  1.20 2.02 1.36 3.48 ;
        RECT  0.10 2.02 0.38 2.30 ;
        RECT  0.16 2.02 0.32 3.48 ;
        END
    END VDD!
    PIN GND!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.00 -0.28 4.80 0.28 ;
        RECT  4.34 -0.28 4.62 0.32 ;
        RECT  3.70 0.68 3.98 0.96 ;
        RECT  3.76 -0.28 3.92 0.96 ;
        RECT  1.16 0.96 1.44 1.24 ;
        RECT  1.22 -0.28 1.38 1.24 ;
        END
    END GND!
    OBS
        LAYER ME1 ;
        RECT  0.10 0.44 0.38 0.72 ;
        RECT  0.22 0.44 0.38 1.24 ;
        RECT  0.22 0.96 0.52 1.24 ;
        RECT  0.22 1.08 0.70 1.24 ;
        RECT  0.54 1.08 0.70 2.30 ;
        RECT  0.54 2.02 0.90 2.30 ;
        RECT  2.08 0.96 2.36 1.24 ;
        RECT  1.78 1.08 2.70 1.24 ;
        RECT  2.54 1.08 2.70 1.74 ;
        RECT  2.54 1.46 2.94 1.74 ;
        RECT  1.78 1.08 1.94 2.30 ;
        RECT  1.66 2.02 1.94 2.30 ;
        RECT  2.86 0.68 3.26 0.96 ;
        RECT  3.10 1.52 4.25 1.68 ;
        RECT  3.97 1.46 4.25 1.74 ;
        RECT  3.10 0.68 3.26 2.25 ;
        RECT  3.10 1.97 3.46 2.25 ;
    END
END AND22NOR2SP1V1_0

END LIBRARY

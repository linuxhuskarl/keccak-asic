/techfiles_ldap/umc_ksmi_lab/techLEF/tech8m2t/tech8m2t.lef
VERSION 5.5 ;

NAMESCASESENSITIVE ON ;

UNITS
    DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID    0.010000 ;

LAYER PO1
    TYPE MASTERSLICE ;
END PO1

LAYER CONT
    TYPE CUT ;
    DCCURRENTDENSITY AVERAGE 0.61 ;
END CONT

LAYER ME1
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;    
    PITCH 0.40 ;
    WIDTH 0.16 ;
    OFFSET 0.0 ;
    AREA 0.1024 ;    
    SPACING 0.16 ;
    SPACING 0.26 RANGE 1.76 1000 ;
    MINIMUMCUT 2 WIDTH 1.4 FROMABOVE ;
    MAXWIDTH 25.0 ;
    MINWIDTH 0.16 ;
    MINENCLOSEDAREA 0.3072 ;
    RESISTANCE RPERSQ 0.0700000000 ;
    CAPACITANCE CPERSQDIST 0.001047 ;
    HEIGHT 0.81 ;
    THICKNESS 0.29 ;
    MINIMUMDENSITY 20.0 ;
    MAXIMUMDENSITY 80.0 ;
    DENSITYCHECKWINDOW 200.0 200.0 ;
    DENSITYCHECKSTEP 100.0 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 400.0 ;
    ANTENNACUMAREARATIO 400.0 ;
    ANTENNAAREAFACTOR 1.0 ;
    ACCURRENTDENSITY RMS 
	FREQUENCY 1 ;
	WIDTH 0.16 ;
	TABLEENTRIES 3.44 ;
    DCCURRENTDENSITY AVERAGE 2.56 ;
END ME1

LAYER VI1
    TYPE CUT ;
    SPACING 0.20 ;
    DCCURRENTDENSITY AVERAGE 0.76 ;
END VI1

LAYER ME2
    TYPE ROUTING ;
    DIRECTION VERTICAL ;
    PITCH 0.40 ;
    WIDTH 0.20 ;
    OFFSET 0.20 ;
    AREA 0.1024 ;
    SPACING 0.20 ;
    SPACING 0.28 RANGE 2 1000 ;
    MINIMUMCUT 2 WIDTH 1.4 ;
    MAXWIDTH 25.0 ;
    MINWIDTH 0.2 ;
    MINENCLOSEDAREA 0.3072 ;
    RESISTANCE RPERSQ 0.0700000000 ;
    CAPACITANCE CPERSQDIST 0.000913 ;
    HEIGHT 14.9 ;
    THICKNESS 0.32 ;
    MINIMUMDENSITY 20.0 ;
    MAXIMUMDENSITY 80.0 ;
    DENSITYCHECKWINDOW 200.0 200.0 ;
    DENSITYCHECKSTEP 100.0 ;
    ANTENNAAREARATIO 400.0 ;
    ANTENNACUMAREARATIO 400.0 ;
    ANTENNAAREAFACTOR 1.0 ;
    ACCURRENTDENSITY RMS 
	FREQUENCY 1 ;
	WIDTH 0.2 ;
	TABLEENTRIES 2.69 ;
    DCCURRENTDENSITY AVERAGE 2.56 ;
END ME2

LAYER VI2
    TYPE CUT ;
    SPACING 0.20 ;
    DCCURRENTDENSITY AVERAGE 0.76 ;
END VI2

LAYER ME3
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;
    PITCH 0.40 ;
    WIDTH 0.20 ;
    OFFSET 0.0 ;
    AREA 0.1024 ;
    SPACING 0.2 ;
    SPACING 0.28 RANGE 2 1000 ;
    MINIMUMCUT 2 WIDTH 1.4 ;
    MAXWIDTH 25.0 ;
    MINWIDTH 0.2 ;
    MINENCLOSEDAREA 0.3072 ;
    RESISTANCE RPERSQ 0.0700000000 ;
    CAPACITANCE CPERSQDIST 0.000912 ;
    HEIGHT 21.7 ;
    THICKNESS 0.32 ;
    MINIMUMDENSITY 20.0 ;
    MAXIMUMDENSITY 80.0 ;
    DENSITYCHECKWINDOW 200.0 200.0 ;
    DENSITYCHECKSTEP 100.0 ;
    ANTENNAAREARATIO 400.0 ;
    ANTENNACUMAREARATIO 400.0 ;
    ANTENNAAREAFACTOR 1.0 ;
    ACCURRENTDENSITY RMS 
	FREQUENCY 1 ;
	WIDTH 0.2 ;
	TABLEENTRIES 2.69 ;
    DCCURRENTDENSITY AVERAGE 2.56 ;
END ME3

LAYER VI3
    TYPE CUT ;
    SPACING 0.20 ;
    DCCURRENTDENSITY AVERAGE 0.76 ;
END VI3

LAYER ME4
    TYPE ROUTING ;
    DIRECTION VERTICAL ;
    PITCH 0.40 ;
    WIDTH 0.20 ;
    OFFSET 0.20 ;
    AREA 0.1024 ;
    SPACING 0.20 ;
    SPACING 0.28 RANGE 2 1000 ;
    MINIMUMCUT 2 WIDTH 1.40 ;
    MAXWIDTH 25.0 ;
    MINWIDTH 0.20 ;
    MINENCLOSEDAREA 0.3072 ;
    RESISTANCE RPERSQ 0.0700000000 ;
    CAPACITANCE CPERSQDIST 0.000914 ;
    HEIGHT 28.5 ;
    THICKNESS 0.32 ;
    MINIMUMDENSITY 20.0 ;
    MAXIMUMDENSITY 80.0 ;
    DENSITYCHECKWINDOW 200.0 200.0 ;
    DENSITYCHECKSTEP 100.0 ;
    ANTENNAAREARATIO 400.0 ;
    ANTENNACUMAREARATIO 400.0 ;
    ANTENNAAREAFACTOR 1.0 ;
    ACCURRENTDENSITY RMS 
	FREQUENCY 1 ;
	WIDTH 0.2 ;
	TABLEENTRIES 2.69 ;
    DCCURRENTDENSITY AVERAGE 2.56 ;
END ME4

LAYER VI4
    TYPE CUT ;
    SPACING 0.20 ;
    DCCURRENTDENSITY AVERAGE 0.76 ;
END VI4

LAYER ME5
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;
    PITCH 0.40 ;
    WIDTH 0.20 ;
    OFFSET 0.0 ;
    AREA 0.1024 ;
    SPACING 0.20 ;
    SPACING 0.28 RANGE 2 1000 ;
    MINIMUMCUT 2 WIDTH 1.40 ;
    MAXWIDTH 25.0 ;
    MINWIDTH 0.20 ;
    MINENCLOSEDAREA 0.3072 ;
    RESISTANCE RPERSQ 0.0700000000 ;
    CAPACITANCE CPERSQDIST 0.000912 ;
    HEIGHT 35.3 ;
    THICKNESS 0.32 ;
    MINIMUMDENSITY 20.0 ;
    MAXIMUMDENSITY 80.0 ;
    DENSITYCHECKWINDOW 200.0 200.0 ;
    DENSITYCHECKSTEP 100.0 ;
    ANTENNAAREARATIO 400.0 ;
    ANTENNACUMAREARATIO 400.0 ;
    ANTENNAAREAFACTOR 1.0 ;
    ACCURRENTDENSITY RMS 
	FREQUENCY 1 ;
	WIDTH 0.2 ;
	TABLEENTRIES 2.69 ;
    DCCURRENTDENSITY AVERAGE 2.56 ;
END ME5

LAYER VI5
    TYPE CUT ;
    SPACING 0.20 ;
    DCCURRENTDENSITY AVERAGE 0.76 ;
END VI5

LAYER ME6
    TYPE ROUTING ;
    DIRECTION VERTICAL ;
    PITCH 0.40 ;
    WIDTH 0.20 ;
    OFFSET 0.20 ;
    AREA 0.1024 ;
    SPACING 0.20 ;
    SPACING 0.28 RANGE 2 1000 ;
    MINIMUMCUT 2 WIDTH 1.40 ;
    MAXWIDTH 25.0 ;
    MINWIDTH 0.20 ;
    MINENCLOSEDAREA 0.3072 ;
    RESISTANCE RPERSQ 0.0700000000 ;
    CAPACITANCE CPERSQDIST 0.000914 ;
    HEIGHT 42.1 ;
    THICKNESS 0.32 ;
    MINIMUMDENSITY 20.0 ;
    MAXIMUMDENSITY 80.0 ;
    DENSITYCHECKWINDOW 200.0 200.0 ;
    DENSITYCHECKSTEP 100.0 ;
    ANTENNAAREARATIO 400.0 ;
    ANTENNACUMAREARATIO 400.0 ;
    ANTENNAAREAFACTOR 1.0 ;
    ACCURRENTDENSITY RMS 
	FREQUENCY 1 ;
	WIDTH 0.2 ;
	TABLEENTRIES 2.69 ;
    DCCURRENTDENSITY AVERAGE 2.56 ;
END ME6

LAYER VI6
    TYPE CUT ;
    SPACING 0.40 ;
    DCCURRENTDENSITY AVERAGE 1.80 ;
END VI6

LAYER ME7
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;
    PITCH 0.80 ;
    WIDTH 0.40 ;
    OFFSET 0.0 ;
    AREA 0.33 ;
    SPACING 0.40 ;
    SPACING 0.5 RANGE 1.60 1000 ;
    MAXWIDTH 25.0 ;
    MINWIDTH 0.40 ;
    MINENCLOSEDAREA 0.87 ;
    RESISTANCE RPERSQ 0.0270000000 ;
    CAPACITANCE CPERSQDIST 0.00052 ;
    HEIGHT 51.45 ;
    THICKNESS 0.8 ;
    MINIMUMDENSITY 20.0 ;
    MAXIMUMDENSITY 80.0 ;
    DENSITYCHECKWINDOW 200.0 200.0 ;
    DENSITYCHECKSTEP 100.0 ;
    ANTENNAAREARATIO 400.0 ;
    ANTENNACUMAREARATIO 400.0 ;
    ANTENNAAREAFACTOR 1.1 ;
    ACCURRENTDENSITY RMS 
	FREQUENCY 1 ;
	WIDTH 0.2 ;
	TABLEENTRIES 6.76 ;
    DCCURRENTDENSITY AVERAGE 8.0 ;
END ME7

LAYER VI7
    TYPE CUT ;
    SPACING 0.40 ;
    DCCURRENTDENSITY AVERAGE 3.60 ;
END VI7

LAYER ME8
    TYPE ROUTING ;
    DIRECTION VERTICAL ;
    PITCH 0.80 ;
    WIDTH 0.40 ;
    OFFSET 0.40 ;
    AREA 0.33 ;
    SPACING 0.40 ;
    SPACING 0.5 RANGE 1.60 1000 ;
    MAXWIDTH 25.0 ;
    MINWIDTH 0.40 ;
    MINENCLOSEDAREA 0.87 ;
    RESISTANCE RPERSQ 0.0270000000 ;
    CAPACITANCE CPERSQDIST 0.00047 ;
    HEIGHT 65.6 ;
    THICKNESS 0.8 ;
    MINIMUMDENSITY 20.0 ;
    MAXIMUMDENSITY 80.0 ;
    DENSITYCHECKWINDOW 200.0 200.0 ;
    DENSITYCHECKSTEP 100.0 ;
    ANTENNAAREARATIO 400.0 ;
    ANTENNACUMAREARATIO 400.0 ;
    ANTENNAAREAFACTOR 1.1 ;
    ACCURRENTDENSITY RMS 
	FREQUENCY 1 ;
	WIDTH 0.2 ;
	TABLEENTRIES 6.76 ;
    DCCURRENTDENSITY AVERAGE 8.0 ;
END ME8

VIA VIA12_HH DEFAULT
    LAYER ME1 ;
        RECT -0.16 -0.10 0.16 0.10 ;
    LAYER VI1 ;
        RECT -0.10 -0.10 0.10 0.10 ;
    LAYER ME2 ;
        RECT -0.16 -0.10 0.16 0.10 ;
    RESISTANCE 1.5 ;
END VIA12_HH

VIA VIA12_HV DEFAULT
    LAYER ME1 ;
        RECT -0.10 -0.16 0.10 0.16 ;
    LAYER VI1 ;
        RECT -0.10 -0.10 0.10 0.10 ;
    LAYER ME2 ;
        RECT -0.16 -0.10 0.16 0.10 ;
    RESISTANCE 1.5 ;
END VIA12_HV

VIA VIA12_VH DEFAULT
    LAYER ME1 ;
        RECT -0.16 -0.10 0.16 0.10 ;
    LAYER VI1 ;
        RECT -0.10 -0.10 0.10 0.10 ;
    LAYER ME2 ;
        RECT -0.10 -0.16 0.10 0.16 ;
    RESISTANCE 1.5 ;
END VIA12_VH

VIA VIA12_VV DEFAULT
    LAYER ME1 ;
        RECT -0.10 -0.16 0.10 0.16 ;
    LAYER VI1 ;
        RECT -0.10 -0.10 0.10 0.10 ;
    LAYER ME2 ;
        RECT -0.10 -0.16 0.10 0.16 ;
    RESISTANCE 1.5 ;
END VIA12_VV

VIA VIA23_HH DEFAULT
    LAYER ME2 ;
        RECT -0.16 -0.10 0.16 0.10 ;
    LAYER VI2 ;
        RECT -0.10 -0.10 0.10 0.10 ;
    LAYER ME3 ;
        RECT -0.16 -0.10 0.16 0.10 ;
    RESISTANCE 1.5 ;
END VIA23_HH

VIA VIA23_HV DEFAULT
    LAYER ME2 ;
        RECT -0.16 -0.10 0.16 0.10 ;
    LAYER VI2 ;
        RECT -0.10 -0.10 0.10 0.10 ;
    LAYER ME3 ;
        RECT -0.10 -0.16 0.10 0.16 ;
    RESISTANCE 1.5 ;
END VIA23_HV

VIA VIA23_VH DEFAULT
    LAYER ME2 ;
        RECT -0.10 -0.16 0.10 0.16 ;
    LAYER VI2 ;
        RECT -0.10 -0.10 0.10 0.10 ;
    LAYER ME3 ;
        RECT -0.16 -0.10 0.16 0.10 ;
    RESISTANCE 1.5 ;
END VIA23_VH

VIA VIA23_VV DEFAULT
    LAYER ME2 ;
        RECT -0.10 -0.16 0.10 0.16 ;
    LAYER VI2 ;
        RECT -0.10 -0.10 0.10 0.10 ;
    LAYER ME3 ;
        RECT -0.10 -0.16 0.10 0.16 ;
    RESISTANCE 1.5 ;
END VIA23_VV

VIA VIA34_HH DEFAULT
    LAYER ME3 ;
        RECT -0.16 -0.10 0.16 0.10 ;
    LAYER VI3 ;
        RECT -0.10 -0.10 0.10 0.10 ;
    LAYER ME4 ;
        RECT -0.16 -0.10 0.16 0.10 ;
    RESISTANCE 1.5 ;
END VIA34_HH

VIA VIA34_HV DEFAULT
    LAYER ME3 ;
        RECT -0.10 -0.16 0.10 0.16 ;
    LAYER VI3 ;
        RECT -0.10 -0.10 0.10 0.10 ;
    LAYER ME4 ;
        RECT -0.16 -0.10 0.16 0.10 ;
    RESISTANCE 1.5 ;
END VIA34_HV

VIA VIA34_VH DEFAULT
    LAYER ME3 ;
        RECT -0.16 -0.10 0.16 0.10 ;
    LAYER VI3 ;
        RECT -0.10 -0.10 0.10 0.10 ;
    LAYER ME4 ;
        RECT -0.10 -0.16 0.10 0.16 ;
    RESISTANCE 1.5 ;
END VIA34_VH

VIA VIA34_VV DEFAULT
    LAYER ME3 ;
        RECT -0.10 -0.16 0.10 0.16 ;
    LAYER VI3 ;
        RECT -0.10 -0.10 0.10 0.10 ;
    LAYER ME4 ;
        RECT -0.10 -0.16 0.10 0.16 ;
    RESISTANCE 1.5 ;
END VIA34_VV

VIA VIA45_HH DEFAULT
    LAYER ME4 ;
        RECT -0.16 -0.10 0.16 0.10 ;
    LAYER VI4 ;
        RECT -0.10 -0.10 0.10 0.10 ;
    LAYER ME5 ;
        RECT -0.16 -0.10 0.16 0.10 ;
    RESISTANCE 1.5 ;
END VIA45_HH

VIA VIA45_HV DEFAULT
    LAYER ME4 ;
        RECT -0.16 -0.10 0.16 0.10 ;
    LAYER VI4 ;
        RECT -0.10 -0.10 0.10 0.10 ;
    LAYER ME5 ;
        RECT -0.10 -0.16 0.10 0.16 ;
    RESISTANCE 1.5 ;
END VIA45_HV

VIA VIA45_VH DEFAULT
    LAYER ME4 ;
        RECT -0.10 -0.16 0.10 0.16 ;
    LAYER VI4 ;
        RECT -0.10 -0.10 0.10 0.10 ;
    LAYER ME5 ;
        RECT -0.16 -0.10 0.16 0.10 ;
    RESISTANCE 1.5 ;
END VIA45_VH

VIA VIA45_VV DEFAULT
    LAYER ME4 ;
        RECT -0.10 -0.16 0.10 0.16 ;
    LAYER VI4 ;
        RECT -0.10 -0.10 0.10 0.10 ;
    LAYER ME5 ;
        RECT -0.10 -0.16 0.10 0.16 ;
    RESISTANCE 1.5 ;
END VIA45_VV

VIA VIA56_HH DEFAULT
    LAYER ME5 ;
        RECT -0.16 -0.10 0.16 0.10 ;
    LAYER VI5 ;
        RECT -0.10 -0.10 0.10 0.10 ;
    LAYER ME6 ;
        RECT -0.16 -0.10 0.16 0.10 ;
    RESISTANCE 1.5 ;
END VIA56_HH

VIA VIA56_HV DEFAULT
    LAYER ME5 ;
        RECT -0.10 -0.16 0.10 0.16 ;
    LAYER VI5 ;
        RECT -0.10 -0.10 0.10 0.10 ;
    LAYER ME6 ;
        RECT -0.16 -0.10 0.16 0.10 ;
    RESISTANCE 1.5 ;
END VIA56_HV

VIA VIA56_VH DEFAULT
    LAYER ME5 ;
        RECT -0.16 -0.10 0.16 0.10 ;
    LAYER VI5 ;
        RECT -0.10 -0.10 0.10 0.10 ;
    LAYER ME6 ;
        RECT -0.10 -0.16 0.10 0.16 ;
    RESISTANCE 1.5 ;
END VIA56_VH

VIA VIA56_VV DEFAULT
    LAYER ME5 ;
        RECT -0.10 -0.16 0.10 0.16 ;
    LAYER VI5 ;
        RECT -0.10 -0.10 0.10 0.10 ;
    LAYER ME6 ;
        RECT -0.10 -0.16 0.10 0.16 ;
    RESISTANCE 1.5 ;
END VIA56_VV

VIA VIA67_DEF DEFAULT
    LAYER ME6 ;
        RECT -0.20 -0.20 0.20 0.20 ;
    LAYER VI6 ;
        RECT -0.20 -0.20 0.20 0.20 ;
    LAYER ME7 ;
        RECT -0.20 -0.20 0.20 0.20 ;
    RESISTANCE 0.6 ;
END VIA67_DEF

VIA VIA78_DEF DEFAULT
    LAYER ME7 ;
        RECT -0.20 -0.20 0.20 0.20 ;
    LAYER VI7 ;
        RECT -0.20 -0.20 0.20 0.20 ;
    LAYER ME8 ;
        RECT -0.20 -0.20 0.20 0.20 ;
    RESISTANCE 0.6 ;
END VIA78_DEF

VIA VIA23_STACK_HAMMER1 DEFAULT TOPOFSTACKONLY
    LAYER ME2 ;
        RECT -0.10 -0.36 0.10 0.16 ;
    LAYER VI2 ;
        RECT -0.10 -0.10 0.10 0.10 ;
    LAYER ME3 ;
        RECT -0.16 -0.10 0.16 0.10 ;
    RESISTANCE 1.5 ;
END VIA23_STACK_HAMMER1

VIA VIA23_STACK_HAMMER2 DEFAULT TOPOFSTACKONLY
    LAYER ME2 ;
        RECT -0.10 -0.16 0.10 0.36 ;
    LAYER VI2 ;
        RECT -0.10 -0.10 0.10 0.10 ;
    LAYER ME3 ;
        RECT -0.16 -0.10 0.16 0.10 ;
    RESISTANCE 1.5 ;
END VIA23_STACK_HAMMER2

VIA VIA23_STACK_CROSS DEFAULT TOPOFSTACKONLY
    LAYER ME2 ;
        RECT -0.10 -0.26 0.10 0.26 ;
    LAYER VI2 ;
        RECT -0.10 -0.10 0.10 0.10 ;
    LAYER ME3 ;
        RECT -0.16 -0.10 0.16 0.10 ;
    RESISTANCE 1.5 ;
END VIA23_STACK_CROSS

VIA VIA34_STACK_HAMMER1 DEFAULT TOPOFSTACKONLY
    LAYER ME3 ;
        RECT -0.36 -0.10 0.16 0.10 ;
    LAYER VI3 ;
        RECT -0.10 -0.10 0.10 0.10 ;
    LAYER ME4 ;
        RECT -0.10 -0.16 0.10 0.16 ;
    RESISTANCE 1.5 ;
END VIA34_STACK_HAMMER1

VIA VIA34_STACK_HAMMER2 DEFAULT TOPOFSTACKONLY
    LAYER ME3 ;
        RECT -0.16 -0.10 0.36 0.10 ;
    LAYER VI3 ;
        RECT -0.10 -0.10 0.10 0.10 ;
    LAYER ME4 ;
        RECT -0.10 -0.16 0.10 0.16 ;
    RESISTANCE 1.5 ;
END VIA34_STACK_HAMMER2

VIA VIA34_STACK_CROSS DEFAULT TOPOFSTACKONLY
    LAYER ME3 ;
        RECT -0.26 -0.10 0.26 0.10 ;
    LAYER VI3 ;
        RECT -0.10 -0.10 0.10 0.10 ;
    LAYER ME4 ;
        RECT -0.10 -0.16 0.10 0.16 ;
    RESISTANCE 1.5 ;
END VIA34_STACK_CROSS

VIA VIA45_STACK_HAMMER1 DEFAULT TOPOFSTACKONLY
    LAYER ME4 ;
        RECT -0.10 -0.36 0.10 0.16 ;
    LAYER VI4 ;
        RECT -0.10 -0.10 0.10 0.10 ;
    LAYER ME5 ;
        RECT -0.16 -0.10 0.16 0.10 ;
    RESISTANCE 1.5 ;
END VIA45_STACK_HAMMER1

VIA VIA45_STACK_HAMMER2 DEFAULT TOPOFSTACKONLY
    LAYER ME4 ;
        RECT -0.10 -0.16 0.10 0.36 ;
    LAYER VI4 ;
        RECT -0.10 -0.10 0.10 0.10 ;
    LAYER ME5 ;
        RECT -0.16 -0.10 0.16 0.10 ;
    RESISTANCE 1.5 ;
END VIA45_STACK_HAMMER2

VIA VIA45_STACK_CROSS DEFAULT TOPOFSTACKONLY
    LAYER ME4 ;
        RECT -0.10 -0.26 0.10 0.26 ;
    LAYER VI4 ;
        RECT -0.10 -0.10 0.10 0.10 ;
    LAYER ME5 ;
        RECT -0.16 -0.10 0.16 0.10 ;
    RESISTANCE 1.5 ;
END VIA45_STACK_CROSS

VIA VIA56_STACK_HAMMER1 DEFAULT TOPOFSTACKONLY
    LAYER ME5 ;
        RECT -0.36 -0.10 0.16 0.10 ;
    LAYER VI5 ;
        RECT -0.10 -0.10 0.10 0.10 ;
    LAYER ME6 ;
        RECT -0.10 -0.16 0.10 0.16 ;
    RESISTANCE 1.5 ;
END VIA56_STACK_HAMMER1

VIA VIA56_STACK_HAMMER2 DEFAULT TOPOFSTACKONLY
    LAYER ME5 ;
        RECT -0.16 -0.10 0.36 0.10 ;
    LAYER VI5 ;
        RECT -0.10 -0.10 0.10 0.10 ;
    LAYER ME6 ;
        RECT -0.10 -0.16 0.10 0.16 ;
    RESISTANCE 1.5 ;
END VIA56_STACK_HAMMER2

VIA VIA56_STACK_CROSS DEFAULT TOPOFSTACKONLY
    LAYER ME5 ;
        RECT -0.26 -0.10 0.26 0.10 ;
    LAYER VI5 ;
        RECT -0.10 -0.10 0.10 0.10 ;
    LAYER ME6 ;
        RECT -0.10 -0.16 0.10 0.16 ;
    RESISTANCE 1.5 ;
END VIA56_STACK_CROSS

VIA VIA67_STACK_DEF DEFAULT TOPOFSTACKONLY
    LAYER ME6 ;
        RECT -0.20 -0.20 0.20 0.20 ;
    LAYER VI6 ;
        RECT -0.20 -0.20 0.20 0.20 ;
    LAYER ME7 ;
        RECT -0.20 -0.20 0.20 0.20 ;
    RESISTANCE 0.6 ;
END VIA67_STACK_DEF

VIA VIA78_STACK_HAMMER1 DEFAULT TOPOFSTACKONLY
    LAYER ME7 ;
        RECT -0.63 -0.20 0.20 0.20 ;
    LAYER VI7 ;
        RECT -0.20 -0.20 0.20 0.20 ;
    LAYER ME8 ;
        RECT -0.20 -0.20 0.20 0.20 ;
    RESISTANCE 0.6 ;
END VIA78_STACK_HAMMER1

VIA VIA78_STACK_HAMMER2 DEFAULT TOPOFSTACKONLY
    LAYER ME7 ;
        RECT -0.20 -0.20 0.63 0.20 ;
    LAYER VI7 ;
        RECT -0.20 -0.20 0.20 0.20 ;
    LAYER ME8 ;
        RECT -0.20 -0.20 0.20 0.20 ;
    RESISTANCE 0.6 ;
END VIA78_STACK_HAMMER2

VIA VIA78_STACK_CROSS DEFAULT TOPOFSTACKONLY
    LAYER ME7 ;
        RECT -0.42 -0.20 0.41 0.20 ;
    LAYER VI7 ;
        RECT -0.20 -0.20 0.20 0.20 ;
    LAYER ME8 ;
        RECT -0.20 -0.20 0.20 0.20 ;
    RESISTANCE 0.6 ;
END VIA78_STACK_CROSS

VIA VIA12_DC_RIGHT DEFAULT
    LAYER ME1 ;
        RECT -0.16 -0.10 0.56 0.10 ;
    LAYER VI1 ;
        RECT 0.30 -0.10 0.50 0.10 ;
        RECT -0.10 -0.10 0.10 0.10 ;
    LAYER ME2 ;
        RECT -0.10 -0.16 0.50 0.16 ;
END VIA12_DC_RIGHT

VIA VIA12_DC_LEFT DEFAULT
    LAYER ME1 ;
        RECT -0.56 -0.10 0.16 0.10 ;
    LAYER VI1 ;
        RECT -0.10 -0.10 0.10 0.10 ;
        RECT -0.50 -0.10 -0.30 0.10 ;
    LAYER ME2 ;
        RECT -0.50 -0.16 0.10 0.16 ;
END VIA12_DC_LEFT

VIA VIA12_DC_TOP DEFAULT
    LAYER ME1 ;
        RECT -0.16 -0.10 0.16 0.50 ;
    LAYER VI1 ;
        RECT -0.10 0.30 0.10 0.50 ;
        RECT -0.10 -0.10 0.10 0.10 ;
    LAYER ME2 ;
        RECT -0.10 -0.16 0.10 0.56 ;
END VIA12_DC_TOP

VIA VIA12_DC_DOWN DEFAULT
    LAYER ME1 ;
        RECT -0.16 -0.50 0.16 0.10 ;
    LAYER VI1 ;
        RECT -0.10 -0.10 0.10 0.10 ;
        RECT -0.10 -0.50 0.10 -0.30 ;
    LAYER ME2 ;
        RECT -0.10 -0.56 0.10 0.16 ;
END VIA12_DC_DOWN

VIA VIA23_DC_RIGHT DEFAULT
    LAYER ME2 ;
        RECT -0.10 -0.16 0.50 0.16 ;
    LAYER VI2 ;
        RECT 0.30 -0.10 0.50 0.10 ;
        RECT -0.10 -0.10 0.10 0.10 ;
    LAYER ME3 ;
        RECT -0.16 -0.10 0.56 0.10 ;
END VIA23_DC_RIGHT

VIA VIA23_DC_LEFT DEFAULT
    LAYER ME2 ;
        RECT -0.50 -0.16 0.10 0.16 ;
    LAYER VI2 ;
        RECT -0.10 -0.10 0.10 0.10 ;
        RECT -0.50 -0.10 -0.30 0.10 ;
    LAYER ME3 ;
        RECT -0.56 -0.10 0.16 0.10 ;
END VIA23_DC_LEFT

VIA VIA23_DC_TOP DEFAULT
    LAYER ME2 ;
        RECT -0.10 -0.16 0.10 0.56 ;
    LAYER VI2 ;
        RECT -0.10 0.30 0.10 0.50 ;
        RECT -0.10 -0.10 0.10 0.10 ;
    LAYER ME3 ;
        RECT -0.16 -0.10 0.16 0.50 ;
END VIA23_DC_TOP

VIA VIA23_DC_DOWN DEFAULT
    LAYER ME2 ;
        RECT -0.10 -0.56 0.10 0.16 ;
    LAYER VI2 ;
        RECT -0.10 -0.10 0.10 0.10 ;
        RECT -0.10 -0.50 0.10 -0.30 ;
    LAYER ME3 ;
        RECT -0.16 -0.50 0.16 0.10 ;
END VIA23_DC_DOWN

VIA VIA34_DC_RIGHT DEFAULT
    LAYER ME3 ;
        RECT -0.16 -0.10 0.56 0.10 ;
    LAYER VI3 ;
        RECT 0.30 -0.10 0.50 0.10 ;
        RECT -0.10 -0.10 0.10 0.10 ;
    LAYER ME4 ;
        RECT -0.10 -0.16 0.50 0.16 ;
END VIA34_DC_RIGHT

VIA VIA34_DC_LEFT DEFAULT
    LAYER ME3 ;
        RECT -0.56 -0.10 0.16 0.10 ;
    LAYER VI3 ;
        RECT -0.10 -0.10 0.10 0.10 ;
        RECT -0.50 -0.10 -0.30 0.10 ;
    LAYER ME4 ;
        RECT -0.50 -0.16 0.10 0.16 ;
END VIA34_DC_LEFT

VIA VIA34_DC_TOP DEFAULT
    LAYER ME3 ;
        RECT -0.16 -0.10 0.16 0.50 ;
    LAYER VI3 ;
        RECT -0.10 0.30 0.10 0.50 ;
        RECT -0.10 -0.10 0.10 0.10 ;
    LAYER ME4 ;
        RECT -0.10 -0.16 0.10 0.56 ;
END VIA34_DC_TOP

VIA VIA34_DC_DOWN DEFAULT
    LAYER ME3 ;
        RECT -0.16 -0.50 0.16 0.10 ;
    LAYER VI3 ;
        RECT -0.10 -0.10 0.10 0.10 ;
        RECT -0.10 -0.50 0.10 -0.30 ;
    LAYER ME4 ;
        RECT -0.10 -0.56 0.10 0.16 ;
END VIA34_DC_DOWN

VIA VIA45_DC_RIGHT DEFAULT
    LAYER ME4 ;
        RECT -0.10 -0.16 0.50 0.16 ;
    LAYER VI4 ;
        RECT 0.30 -0.10 0.50 0.10 ;
        RECT -0.10 -0.10 0.10 0.10 ;
    LAYER ME5 ;
        RECT -0.16 -0.10 0.56 0.10 ;
END VIA45_DC_RIGHT

VIA VIA45_DC_LEFT DEFAULT
    LAYER ME4 ;
        RECT -0.50 -0.16 0.10 0.16 ;
    LAYER VI4 ;
        RECT -0.10 -0.10 0.10 0.10 ;
        RECT -0.50 -0.10 -0.30 0.10 ;
    LAYER ME5 ;
        RECT -0.56 -0.10 0.16 0.10 ;
END VIA45_DC_LEFT

VIA VIA45_DC_TOP DEFAULT
    LAYER ME4 ;
        RECT -0.10 -0.16 0.10 0.56 ;
    LAYER VI4 ;
        RECT -0.10 0.30 0.10 0.50 ;
        RECT -0.10 -0.10 0.10 0.10 ;
    LAYER ME5 ;
        RECT -0.16 -0.10 0.16 0.50 ;
END VIA45_DC_TOP

VIA VIA45_DC_DOWN DEFAULT
    LAYER ME4 ;
        RECT -0.10 -0.56 0.10 0.16 ;
    LAYER VI4 ;
        RECT -0.10 -0.10 0.10 0.10 ;
        RECT -0.10 -0.50 0.10 -0.30 ;
    LAYER ME5 ;
        RECT -0.16 -0.50 0.16 0.10 ;
END VIA45_DC_DOWN

VIA VIA56_DC_RIGHT DEFAULT
    LAYER ME5 ;
        RECT -0.10 -0.16 0.50 0.16 ;
    LAYER VI5 ;
        RECT 0.30 -0.10 0.50 0.10 ;
        RECT -0.10 -0.10 0.10 0.10 ;
    LAYER ME6 ;
        RECT -0.16 -0.10 0.56 0.10 ;
END VIA56_DC_RIGHT

VIA VIA56_DC_LEFT DEFAULT
    LAYER ME5 ;
        RECT -0.50 -0.16 0.10 0.16 ;
    LAYER VI5 ;
        RECT -0.10 -0.10 0.10 0.10 ;
        RECT -0.50 -0.10 -0.30 0.10 ;
    LAYER ME6 ;
        RECT -0.56 -0.10 0.16 0.10 ;
END VIA56_DC_LEFT

VIA VIA56_DC_TOP DEFAULT
    LAYER ME5 ;
        RECT -0.10 -0.16 0.10 0.56 ;
    LAYER VI5 ;
        RECT -0.10 0.30 0.10 0.50 ;
        RECT -0.10 -0.10 0.10 0.10 ;
    LAYER ME6 ;
        RECT -0.16 -0.10 0.16 0.50 ;
END VIA56_DC_TOP

VIA VIA56_DC_DOWN DEFAULT
    LAYER ME5 ;
        RECT -0.10 -0.56 0.10 0.16 ;
    LAYER VI5 ;
        RECT -0.10 -0.10 0.10 0.10 ;
        RECT -0.10 -0.50 0.10 -0.30 ;
    LAYER ME6 ;
        RECT -0.16 -0.50 0.16 0.10 ;
END VIA56_DC_DOWN

VIA VIA67_DC_RIGHT DEFAULT
    LAYER ME6 ;
        RECT -0.20 -0.20 1.00 0.20 ;
    LAYER VI6 ;
        RECT 0.60 -0.20 1.00 0.20 ;
        RECT -0.20 -0.20 0.20 0.20 ;
    LAYER ME7 ;
        RECT -0.20 -0.20 1.00 0.20 ;
END VIA67_DC_RIGHT

VIA VIA67_DC_LEFT DEFAULT
    LAYER ME6 ;
        RECT -1.00 -0.20 0.20 0.20 ;
    LAYER VI6 ;
        RECT -0.20 -0.20 0.20 0.20 ;
        RECT -1.00 -0.20 -0.60 0.20 ;
    LAYER ME7 ;
        RECT -1.00 -0.20 0.20 0.20 ;
END VIA67_DC_LEFT

VIA VIA67_DC_TOP DEFAULT
    LAYER ME6 ;
        RECT -0.20 -0.20 0.20 1.00 ;
    LAYER VI6 ;
        RECT -0.20 0.60 0.20 1.00 ;
        RECT -0.20 -0.20 0.20 0.20 ;
    LAYER ME7 ;
        RECT -0.20 -0.20 0.20 1.00 ;
END VIA67_DC_TOP

VIA VIA67_DC_DOWN DEFAULT
    LAYER ME6 ;
        RECT -0.20 -1.00 0.20 0.20 ;
    LAYER VI6 ;
        RECT -0.20 -0.20 0.20 0.20 ;
        RECT -0.20 -1.00 0.20 -0.60 ;
    LAYER ME7 ;
        RECT -0.20 -1.00 0.20 0.20 ;
END VIA67_DC_DOWN

VIA VIA78_DC_RIGHT DEFAULT
    LAYER ME7 ;
        RECT -0.20 -0.20 1.00 0.20 ;
    LAYER VI7 ;
        RECT 0.60 -0.20 1.00 0.20 ;
        RECT -0.20 -0.20 0.20 0.20 ;
    LAYER ME8 ;
        RECT -0.20 -0.20 1.00 0.20 ;
END VIA78_DC_RIGHT

VIA VIA78_DC_LEFT DEFAULT
    LAYER ME7 ;
        RECT -1.00 -0.20 0.20 0.20 ;
    LAYER VI7 ;
        RECT -0.20 -0.20 0.20 0.20 ;
        RECT -1.00 -0.20 -0.60 0.20 ;
    LAYER ME8 ;
        RECT -1.00 -0.20 0.20 0.20 ;
END VIA78_DC_LEFT

VIA VIA78_DC_TOP DEFAULT
    LAYER ME7 ;
        RECT -0.20 -0.20 0.20 1.00 ;
    LAYER VI7 ;
        RECT -0.20 0.60 0.20 1.00 ;
        RECT -0.20 -0.20 0.20 0.20 ;
    LAYER ME8 ;
        RECT -0.20 -0.20 0.20 1.00 ;
END VIA78_DC_TOP

VIA VIA78_DC_DOWN DEFAULT
    LAYER ME7 ;
        RECT -0.20 -1.00 0.20 0.20 ;
    LAYER VI7 ;
        RECT -0.20 -0.20 0.20 0.20 ;
        RECT -0.20 -1.00 0.20 -0.60 ;
    LAYER ME8 ;
        RECT -0.20 -1.00 0.20 0.20 ;
END VIA78_DC_DOWN

SPACING
    SAMENET CONT VI1 0 STACK ;
    SAMENET ME1 ME1 0.160000 STACK ;
    SAMENET VI1 VI1 0.200000  ;
    SAMENET ME2 ME2 0.200000 STACK ;
    SAMENET VI1 VI2 0.000000 STACK ;
    SAMENET VI2 VI2 0.200000  ;
    SAMENET ME3 ME3 0.200000 STACK ;
    SAMENET VI2 VI3 0.000000 STACK ;
    SAMENET VI3 VI3 0.200000  ;
    SAMENET ME4 ME4 0.200000 STACK ;
    SAMENET VI3 VI4 0.000000 STACK ;
    SAMENET VI4 VI4 0.200000  ;
    SAMENET ME5 ME5 0.200000 STACK ;
    SAMENET VI4 VI5 0.000000 STACK ;
    SAMENET VI5 VI5 0.200000  ;
    SAMENET ME6 ME6 0.200000 STACK ;
    SAMENET VI5 VI6 0.000000 STACK ;
    SAMENET VI6 VI6 0.400000  ;
    SAMENET ME7 ME7 0.400000 STACK ;
    SAMENET VI6 VI7 0.000000 STACK ;
    SAMENET VI7 VI7 0.400000  ;
    SAMENET ME8 ME8 0.400000  ;
END SPACING

VIARULE VIAM1M2A
    LAYER ME2 ;
        DIRECTION VERTICAL ;
        WIDTH 0.20 TO 0.20 ;

    LAYER ME1 ;
        DIRECTION HORIZONTAL ;
        WIDTH 0.16 TO 0.16 ;
    VIA VIA12_VH ;
    VIA VIA12_HV ;
    VIA VIA12_VV ;
    VIA VIA12_HH ;
END VIAM1M2A

VIARULE VIAM2M3
    LAYER ME3 ;
        DIRECTION HORIZONTAL ;
        WIDTH 0.20 TO 0.20 ;

    LAYER ME2 ;
        DIRECTION VERTICAL ;
        WIDTH 0.20 TO 0.20 ;
    VIA VIA23_HH ;
    VIA VIA23_VV ;
    VIA VIA23_HV ;
    VIA VIA23_VH ;
END VIAM2M3

VIARULE VIAM3M4
    LAYER ME4 ;
        DIRECTION VERTICAL ;
        WIDTH 0.20 TO 0.20 ;

    LAYER ME3 ;
        DIRECTION HORIZONTAL ;
        WIDTH 0.20 TO 0.20 ;
    VIA VIA34_HH ;
    VIA VIA34_VH ;
    VIA VIA34_HV ;
    VIA VIA34_VV ;
END VIAM3M4

VIARULE VIAM4M5
    LAYER ME5 ;
        DIRECTION HORIZONTAL ;
        WIDTH 0.20 TO 0.20 ;

    LAYER ME4 ;
        DIRECTION VERTICAL ;
        WIDTH 0.20 TO 0.20 ;
    VIA VIA45_HV ;
    VIA VIA45_HH ;
    VIA VIA45_VV ;
    VIA VIA45_VH ;
END VIAM4M5

VIARULE VIAM5M6
    LAYER ME6 ;
        DIRECTION VERTICAL ;
        WIDTH 0.40 TO 0.40 ;

    LAYER ME5 ;
        DIRECTION HORIZONTAL ;
        WIDTH 0.20 TO 0.20 ;
    VIA VIA56_VH ;
    VIA VIA56_VV ;
    VIA VIA56_HH ;
    VIA VIA56_HV ;
END VIAM5M6

VIARULE VIAM6M7
    LAYER ME7 ;
        DIRECTION HORIZONTAL ;
        WIDTH 0.40 TO 0.40 ;

    LAYER ME6 ;
        DIRECTION VERTICAL ;
        WIDTH 0.20 TO 0.20 ;
    VIA VIA67_DEF ;
END VIAM6M7

VIARULE VIAM7M8
    LAYER ME8 ;
        DIRECTION VERTICAL ;
        WIDTH 0.40 TO 0.40 ;

    LAYER ME7 ;
        DIRECTION HORIZONTAL ;
        WIDTH 0.40 TO 0.40 ;
    VIA VIA78_DEF ;
END VIAM7M8

VIARULE TURN1 GENERATE
    LAYER ME1 ;
        DIRECTION HORIZONTAL ;

    LAYER ME1 ;
        DIRECTION VERTICAL ;
END TURN1

VIARULE TURN2 GENERATE
    LAYER ME2 ;
        DIRECTION VERTICAL ;

    LAYER ME2 ;
        DIRECTION HORIZONTAL ;
END TURN2

VIARULE TURN3 GENERATE
    LAYER ME3 ;
        DIRECTION VERTICAL ;

    LAYER ME3 ;
        DIRECTION HORIZONTAL ;
END TURN3

VIARULE TURN4 GENERATE
    LAYER ME4 ;
        DIRECTION VERTICAL ;

    LAYER ME4 ;
        DIRECTION HORIZONTAL ;
END TURN4

VIARULE TURN5 GENERATE
    LAYER ME5 ;
        DIRECTION VERTICAL ;

    LAYER ME5 ;
        DIRECTION HORIZONTAL ;
END TURN5

VIARULE TURN6 GENERATE
    LAYER ME6 ;
        DIRECTION VERTICAL ;

    LAYER ME6 ;
        DIRECTION HORIZONTAL ;
END TURN6

VIARULE TURN7 GENERATE
    LAYER ME7 ;
        DIRECTION VERTICAL ;

    LAYER ME7 ;
        DIRECTION HORIZONTAL ;
END TURN7

VIARULE TURN8 GENERATE
    LAYER ME8 ;
        DIRECTION VERTICAL ;

    LAYER ME8 ;
        DIRECTION HORIZONTAL ;
END TURN8

VIARULE GENM1M2A GENERATE
    LAYER ME2 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.06 ;
        METALOVERHANG 0.00 ;

    LAYER ME1 ;
        DIRECTION HORIZONTAL ;
        WIDTH 0.01 TO 1.11 ;
        OVERHANG 0.06 ;
        METALOVERHANG 0.00 ;

    LAYER VI1 ;
        RECT -0.10 -0.10 0.10 0.10 ;
        SPACING 0.40 BY 0.40 ;
END GENM1M2A

VIARULE GENM1M2B GENERATE
    LAYER ME2 ;
        DIRECTION VERTICAL ;
        WIDTH 0.01 TO 1.11 ;
        OVERHANG 0.06 ;
        METALOVERHANG 0.00 ;

    LAYER ME1 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.06 ;
        METALOVERHANG 0.00 ;

    LAYER VI1 ;
        RECT -0.10 -0.10 0.10 0.10 ;
        SPACING 0.40 BY 0.40 ;
END GENM1M2B

VIARULE GENM2M3A GENERATE
    LAYER ME3 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.06 ;
        METALOVERHANG 0.00 ;

    LAYER ME2 ;
        DIRECTION VERTICAL ;
        WIDTH 0.01 TO 1.11 ;
        OVERHANG 0.06 ;
        METALOVERHANG 0.00 ;

    LAYER VI2 ;
        RECT -0.10 -0.10 0.10 0.10 ;
        SPACING 0.40 BY 0.40 ;
END GENM2M3A

VIARULE GENM2M3B GENERATE
    LAYER ME3 ;
        DIRECTION HORIZONTAL ;
        WIDTH 0.01 TO 1.11 ;
        OVERHANG 0.06 ;
        METALOVERHANG 0.00 ;

    LAYER ME2 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.06 ;
        METALOVERHANG 0.00 ;

    LAYER VI2 ;
        RECT -0.10 -0.10 0.10 0.10 ;
        SPACING 0.40 BY 0.40 ;
END GENM2M3B

VIARULE GENM3M4A GENERATE
    LAYER ME4 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.06 ;
        METALOVERHANG 0.00 ;

    LAYER ME3 ;
        DIRECTION HORIZONTAL ;
        WIDTH 0.01 TO 1.11 ;
        OVERHANG 0.06 ;
        METALOVERHANG 0.00 ;

    LAYER VI3 ;
        RECT -0.10 -0.10 0.10 0.10 ;
        SPACING 0.40 BY 0.40 ;
END GENM3M4A

VIARULE GENM3M4B GENERATE
    LAYER ME4 ;
        DIRECTION VERTICAL ;
        WIDTH 0.01 TO 1.11 ;
        OVERHANG 0.06 ;
        METALOVERHANG 0.00 ;

    LAYER ME3 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.06 ;
        METALOVERHANG 0.00 ;

    LAYER VI3 ;
        RECT -0.10 -0.10 0.10 0.10 ;
        SPACING 0.40 BY 0.40 ;
END GENM3M4B

VIARULE GENM4M5A GENERATE
    LAYER ME5 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.06 ;
        METALOVERHANG 0.00 ;

    LAYER ME4 ;
        DIRECTION VERTICAL ;
        WIDTH 0.01 TO 1.11 ;
        OVERHANG 0.06 ;
        METALOVERHANG 0.00 ;

    LAYER VI4 ;
        RECT -0.10 -0.10 0.10 0.10 ;
        SPACING 0.40 BY 0.40 ;
END GENM4M5A

VIARULE GENM4M5B GENERATE
    LAYER ME5 ;
        DIRECTION HORIZONTAL ;
        WIDTH 0.01 TO 1.11 ;
        OVERHANG 0.06 ;
        METALOVERHANG 0.00 ;

    LAYER ME4 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.06 ;
        METALOVERHANG 0.00 ;

    LAYER VI4 ;
        RECT -0.10 -0.10 0.10 0.10 ;
        SPACING 0.40 BY 0.40 ;
END GENM4M5B

VIARULE GENM5M6A GENERATE
    LAYER ME6 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.06 ;
        METALOVERHANG 0.00 ;

    LAYER ME5 ;
        DIRECTION HORIZONTAL ;
        WIDTH 0.01 TO 1.11 ;
        OVERHANG 0.06 ;
        METALOVERHANG 0.00 ;

    LAYER VI5 ;
        RECT -0.10 -0.10 0.10 0.10 ;
        SPACING 0.40 BY 0.40 ;
END GENM5M6A

VIARULE GENM5M6B GENERATE
    LAYER ME6 ;
        DIRECTION VERTICAL ;
        WIDTH 0.01 TO 1.11 ;
        OVERHANG 0.06 ;
        METALOVERHANG 0.00 ;

    LAYER ME5 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.06 ;
        METALOVERHANG 0.00 ;

    LAYER VI5 ;
        RECT -0.10 -0.10 0.10 0.10 ;
        SPACING 0.40 BY 0.40 ;
END GENM5M6B

VIARULE GENM6M7A GENERATE
    LAYER ME7 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.00 ;
        METALOVERHANG 0.00 ;

    LAYER ME6 ;
        DIRECTION HORIZONTAL ;
        WIDTH 0.01 TO 1.99 ;
        OVERHANG 0.00 ;
        METALOVERHANG 0.00 ;

    LAYER VI6 ;
        RECT -0.20 -0.20 0.20 0.20 ;
        SPACING 0.80 BY 0.80 ;
END GENM6M7A

VIARULE GENM6M7B GENERATE
    LAYER ME7 ;
        DIRECTION VERTICAL ;
        WIDTH 0.01 TO 1.99 ;
        OVERHANG 0.00 ;
        METALOVERHANG 0.00 ;

    LAYER ME6 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.00 ;
        METALOVERHANG 0.00 ;

    LAYER VI6 ;
        RECT -0.20 -0.20 0.20 0.20 ;
        SPACING 0.80 BY 0.80 ;
END GENM6M7B

VIARULE GENM7M8A GENERATE
    LAYER ME8 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.00 ;
        METALOVERHANG 0.00 ;

    LAYER ME7 ;
        DIRECTION HORIZONTAL ;
        WIDTH 0.01 TO 1.99 ;
        OVERHANG 0.00 ;
        METALOVERHANG 0.00 ;

    LAYER VI7 ;
        RECT -0.20 -0.20 0.20 0.20 ;
        SPACING 0.80 BY 0.80 ;
END GENM7M8A

VIARULE GENM7M8B GENERATE
    LAYER ME8 ;
        DIRECTION VERTICAL ;
        WIDTH 0.01 TO 1.99 ;
        OVERHANG 0.00 ;
        METALOVERHANG 0.00 ;

    LAYER ME7 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.00 ;
        METALOVERHANG 0.00 ;

    LAYER VI7 ;
        RECT -0.20 -0.20 0.20 0.20 ;
        SPACING 0.80 BY 0.80 ;
END GENM7M8B

VIARULE GENM1M2_W GENERATE
    LAYER ME2 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.06 ;
        METALOVERHANG 0.00 ;

    LAYER ME1 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.06 ;
        METALOVERHANG 0.00 ;

    LAYER VI1 ;
        RECT -0.10 -0.10 0.10 0.10 ;
        SPACING 0.48 BY 0.48 ;
END GENM1M2_W

VIARULE GENM2M3_W GENERATE
    LAYER ME3 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.06 ;
        METALOVERHANG 0.00 ;

    LAYER ME2 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.06 ;
        METALOVERHANG 0.00 ;

    LAYER VI2 ;
        RECT -0.10 -0.10 0.10 0.10 ;
        SPACING 0.48 BY 0.48 ;
END GENM2M3_W

VIARULE GENM3M4_W GENERATE
    LAYER ME4 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.06 ;
        METALOVERHANG 0.00 ;

    LAYER ME3 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.06 ;
        METALOVERHANG 0.00 ;

    LAYER VI3 ;
        RECT -0.10 -0.10 0.10 0.10 ;
        SPACING 0.48 BY 0.48 ;
END GENM3M4_W

VIARULE GENM4M5_W GENERATE
    LAYER ME5 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.06 ;
        METALOVERHANG 0.00 ;

    LAYER ME4 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.06 ;
        METALOVERHANG 0.00 ;

    LAYER VI4 ;
        RECT -0.10 -0.10 0.10 0.10 ;
        SPACING 0.48 BY 0.48 ;
END GENM4M5_W

VIARULE GENM5M6_W GENERATE
    LAYER ME6 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.06 ;
        METALOVERHANG 0.00 ;

    LAYER ME5 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.06 ;
        METALOVERHANG 0.00 ;

    LAYER VI5 ;
        RECT -0.10 -0.10 0.10 0.10 ;
        SPACING 0.48 BY 0.48 ;
END GENM5M6_W

VIARULE GENM6M7_W GENERATE
    LAYER ME7 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.00 ;
        METALOVERHANG 0.00 ;

    LAYER ME6 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.00 ;
        METALOVERHANG 0.00 ;

    LAYER VI6 ;
        RECT -0.20 -0.20 0.20 0.20 ;
        SPACING 0.90 BY 0.90 ;
END GENM6M7_W

VIARULE GENM7M8_W GENERATE
    LAYER ME8 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.00 ;
        METALOVERHANG 0.00 ;

    LAYER ME7 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.00 ;
        METALOVERHANG 0.00 ;

    LAYER VI7 ;
        RECT -0.20 -0.20 0.20 0.20 ;
        SPACING 0.90 BY 0.90 ;
END GENM7M8_W

SITE CoreSite
    SYMMETRY Y  ;
    CLASS CORE  ;
    SIZE 0.40 BY 3.20 ;
END CoreSite

END LIBRARY

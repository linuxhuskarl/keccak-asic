/techfiles_ldap/umc_ksmi_lab/cellsLEF/cells.lef